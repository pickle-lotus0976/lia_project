module lia_digital_core (adc_valid,
    clk,
    mixer_valid,
    rst_n,
    adc_data,
    mixer_i_out,
    mixer_q_out,
    phase_increment);
 input adc_valid;
 input clk;
 output mixer_valid;
 input rst_n;
 input [11:0] adc_data;
 output [23:0] mixer_i_out;
 output [23:0] mixer_q_out;
 input [31:0] phase_increment;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire clknet_leaf_0_clk;
 wire \mixer_i.adc_reg[0] ;
 wire \mixer_i.adc_reg[10] ;
 wire \mixer_i.adc_reg[11] ;
 wire \mixer_i.adc_reg[1] ;
 wire \mixer_i.adc_reg[2] ;
 wire \mixer_i.adc_reg[3] ;
 wire \mixer_i.adc_reg[4] ;
 wire \mixer_i.adc_reg[5] ;
 wire \mixer_i.adc_reg[6] ;
 wire \mixer_i.adc_reg[7] ;
 wire \mixer_i.adc_reg[8] ;
 wire \mixer_i.adc_reg[9] ;
 wire \mixer_i.nco_data[0] ;
 wire \mixer_i.nco_data[10] ;
 wire \mixer_i.nco_data[11] ;
 wire \mixer_i.nco_data[1] ;
 wire \mixer_i.nco_data[2] ;
 wire \mixer_i.nco_data[3] ;
 wire \mixer_i.nco_data[4] ;
 wire \mixer_i.nco_data[5] ;
 wire \mixer_i.nco_data[6] ;
 wire \mixer_i.nco_data[7] ;
 wire \mixer_i.nco_data[8] ;
 wire \mixer_i.nco_data[9] ;
 wire \mixer_i.nco_reg[0] ;
 wire \mixer_i.nco_reg[10] ;
 wire \mixer_i.nco_reg[11] ;
 wire \mixer_i.nco_reg[1] ;
 wire \mixer_i.nco_reg[2] ;
 wire \mixer_i.nco_reg[3] ;
 wire \mixer_i.nco_reg[4] ;
 wire \mixer_i.nco_reg[5] ;
 wire \mixer_i.nco_reg[6] ;
 wire \mixer_i.nco_reg[7] ;
 wire \mixer_i.nco_reg[8] ;
 wire \mixer_i.nco_reg[9] ;
 wire \mixer_i.nco_valid ;
 wire \mixer_i.product[0] ;
 wire \mixer_i.product[10] ;
 wire \mixer_i.product[11] ;
 wire \mixer_i.product[12] ;
 wire \mixer_i.product[13] ;
 wire \mixer_i.product[14] ;
 wire \mixer_i.product[15] ;
 wire \mixer_i.product[16] ;
 wire \mixer_i.product[17] ;
 wire \mixer_i.product[18] ;
 wire \mixer_i.product[19] ;
 wire \mixer_i.product[1] ;
 wire \mixer_i.product[20] ;
 wire \mixer_i.product[21] ;
 wire \mixer_i.product[22] ;
 wire \mixer_i.product[23] ;
 wire \mixer_i.product[2] ;
 wire \mixer_i.product[3] ;
 wire \mixer_i.product[4] ;
 wire \mixer_i.product[5] ;
 wire \mixer_i.product[6] ;
 wire \mixer_i.product[7] ;
 wire \mixer_i.product[8] ;
 wire \mixer_i.product[9] ;
 wire \mixer_i.product_delayed[0] ;
 wire \mixer_i.product_delayed[10] ;
 wire \mixer_i.product_delayed[11] ;
 wire \mixer_i.product_delayed[12] ;
 wire \mixer_i.product_delayed[13] ;
 wire \mixer_i.product_delayed[14] ;
 wire \mixer_i.product_delayed[15] ;
 wire \mixer_i.product_delayed[16] ;
 wire \mixer_i.product_delayed[17] ;
 wire \mixer_i.product_delayed[18] ;
 wire \mixer_i.product_delayed[19] ;
 wire \mixer_i.product_delayed[1] ;
 wire \mixer_i.product_delayed[20] ;
 wire \mixer_i.product_delayed[21] ;
 wire \mixer_i.product_delayed[22] ;
 wire \mixer_i.product_delayed[23] ;
 wire \mixer_i.product_delayed[2] ;
 wire \mixer_i.product_delayed[3] ;
 wire \mixer_i.product_delayed[4] ;
 wire \mixer_i.product_delayed[5] ;
 wire \mixer_i.product_delayed[6] ;
 wire \mixer_i.product_delayed[7] ;
 wire \mixer_i.product_delayed[8] ;
 wire \mixer_i.product_delayed[9] ;
 wire \mixer_i.valid_stage1 ;
 wire \mixer_i.valid_stage2 ;
 wire \mixer_i.valid_stage2_delayed ;
 wire \mixer_q.nco_data[0] ;
 wire \mixer_q.nco_data[10] ;
 wire \mixer_q.nco_data[11] ;
 wire \mixer_q.nco_data[1] ;
 wire \mixer_q.nco_data[2] ;
 wire \mixer_q.nco_data[3] ;
 wire \mixer_q.nco_data[4] ;
 wire \mixer_q.nco_data[5] ;
 wire \mixer_q.nco_data[6] ;
 wire \mixer_q.nco_data[7] ;
 wire \mixer_q.nco_data[8] ;
 wire \mixer_q.nco_data[9] ;
 wire \mixer_q.nco_reg[0] ;
 wire \mixer_q.nco_reg[10] ;
 wire \mixer_q.nco_reg[11] ;
 wire \mixer_q.nco_reg[1] ;
 wire \mixer_q.nco_reg[2] ;
 wire \mixer_q.nco_reg[3] ;
 wire \mixer_q.nco_reg[4] ;
 wire \mixer_q.nco_reg[5] ;
 wire \mixer_q.nco_reg[6] ;
 wire \mixer_q.nco_reg[7] ;
 wire \mixer_q.nco_reg[8] ;
 wire \mixer_q.nco_reg[9] ;
 wire \mixer_q.product[0] ;
 wire \mixer_q.product[10] ;
 wire \mixer_q.product[11] ;
 wire \mixer_q.product[12] ;
 wire \mixer_q.product[13] ;
 wire \mixer_q.product[14] ;
 wire \mixer_q.product[15] ;
 wire \mixer_q.product[16] ;
 wire \mixer_q.product[17] ;
 wire \mixer_q.product[18] ;
 wire \mixer_q.product[19] ;
 wire \mixer_q.product[1] ;
 wire \mixer_q.product[20] ;
 wire \mixer_q.product[21] ;
 wire \mixer_q.product[22] ;
 wire \mixer_q.product[23] ;
 wire \mixer_q.product[2] ;
 wire \mixer_q.product[3] ;
 wire \mixer_q.product[4] ;
 wire \mixer_q.product[5] ;
 wire \mixer_q.product[6] ;
 wire \mixer_q.product[7] ;
 wire \mixer_q.product[8] ;
 wire \mixer_q.product[9] ;
 wire \mixer_q.product_delayed[0] ;
 wire \mixer_q.product_delayed[10] ;
 wire \mixer_q.product_delayed[11] ;
 wire \mixer_q.product_delayed[12] ;
 wire \mixer_q.product_delayed[13] ;
 wire \mixer_q.product_delayed[14] ;
 wire \mixer_q.product_delayed[15] ;
 wire \mixer_q.product_delayed[16] ;
 wire \mixer_q.product_delayed[17] ;
 wire \mixer_q.product_delayed[18] ;
 wire \mixer_q.product_delayed[19] ;
 wire \mixer_q.product_delayed[1] ;
 wire \mixer_q.product_delayed[20] ;
 wire \mixer_q.product_delayed[21] ;
 wire \mixer_q.product_delayed[22] ;
 wire \mixer_q.product_delayed[23] ;
 wire \mixer_q.product_delayed[2] ;
 wire \mixer_q.product_delayed[3] ;
 wire \mixer_q.product_delayed[4] ;
 wire \mixer_q.product_delayed[5] ;
 wire \mixer_q.product_delayed[6] ;
 wire \mixer_q.product_delayed[7] ;
 wire \mixer_q.product_delayed[8] ;
 wire \mixer_q.product_delayed[9] ;
 wire \nco_inst.cosine_lut.addr[0] ;
 wire \nco_inst.cosine_lut.addr[1] ;
 wire \nco_inst.cosine_lut.addr[2] ;
 wire \nco_inst.cosine_lut.addr[3] ;
 wire \nco_inst.cosine_lut.addr[4] ;
 wire \nco_inst.cosine_lut.addr[5] ;
 wire \nco_inst.lut_addr_sin[6] ;
 wire \nco_inst.lut_addr_sin[7] ;
 wire \nco_inst.phase_accum[0] ;
 wire \nco_inst.phase_accum[10] ;
 wire \nco_inst.phase_accum[11] ;
 wire \nco_inst.phase_accum[12] ;
 wire \nco_inst.phase_accum[13] ;
 wire \nco_inst.phase_accum[14] ;
 wire \nco_inst.phase_accum[15] ;
 wire \nco_inst.phase_accum[16] ;
 wire \nco_inst.phase_accum[17] ;
 wire \nco_inst.phase_accum[18] ;
 wire \nco_inst.phase_accum[19] ;
 wire \nco_inst.phase_accum[1] ;
 wire \nco_inst.phase_accum[20] ;
 wire \nco_inst.phase_accum[21] ;
 wire \nco_inst.phase_accum[22] ;
 wire \nco_inst.phase_accum[23] ;
 wire \nco_inst.phase_accum[2] ;
 wire \nco_inst.phase_accum[3] ;
 wire \nco_inst.phase_accum[4] ;
 wire \nco_inst.phase_accum[5] ;
 wire \nco_inst.phase_accum[6] ;
 wire \nco_inst.phase_accum[7] ;
 wire \nco_inst.phase_accum[8] ;
 wire \nco_inst.phase_accum[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_0_clk;
 wire clknet_2_0_0_clk;
 wire clknet_2_1_0_clk;
 wire clknet_2_2_0_clk;
 wire clknet_2_3_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net904;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net917;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;

 sky130_fd_sc_hd__nand2_1 _3539_ (.A(net257),
    .B(net170),
    .Y(_1147_));
 sky130_fd_sc_hd__buf_2 _3540_ (.A(_1147_),
    .X(_1156_));
 sky130_fd_sc_hd__clkbuf_4 _3541_ (.A(_1156_),
    .X(_1165_));
 sky130_fd_sc_hd__o21ai_1 _3542_ (.A1(net163),
    .A2(net156),
    .B1(net256),
    .Y(_1174_));
 sky130_fd_sc_hd__buf_2 _3543_ (.A(_1174_),
    .X(_1183_));
 sky130_fd_sc_hd__clkbuf_4 _3544_ (.A(_1183_),
    .X(_1193_));
 sky130_fd_sc_hd__nand4_4 _3545_ (.A(net297),
    .B(net284),
    .C(net145),
    .D(net140),
    .Y(_1202_));
 sky130_fd_sc_hd__nand2_1 _3546_ (.A(net273),
    .B(net151),
    .Y(_1212_));
 sky130_fd_sc_hd__nand2_1 _3547_ (.A(net283),
    .B(net145),
    .Y(_1221_));
 sky130_fd_sc_hd__nand2_2 _3548_ (.A(net297),
    .B(net140),
    .Y(_1231_));
 sky130_fd_sc_hd__nand2_2 _3549_ (.A(_1221_),
    .B(_1231_),
    .Y(_1240_));
 sky130_fd_sc_hd__a21boi_2 _3550_ (.A1(_1202_),
    .A2(_1212_),
    .B1_N(_1240_),
    .Y(_1249_));
 sky130_fd_sc_hd__nand2_1 _3551_ (.A(net272),
    .B(net145),
    .Y(_1259_));
 sky130_fd_sc_hd__nand2_1 _3552_ (.A(net283),
    .B(net137),
    .Y(_1268_));
 sky130_fd_sc_hd__nand2_2 _3553_ (.A(_1259_),
    .B(_1268_),
    .Y(_1277_));
 sky130_fd_sc_hd__nand4_1 _3554_ (.A(net283),
    .B(net272),
    .C(net145),
    .D(net138),
    .Y(_1287_));
 sky130_fd_sc_hd__and2_1 _3555_ (.A(net258),
    .B(net151),
    .X(_1296_));
 sky130_fd_sc_hd__a21oi_1 _3556_ (.A1(_1277_),
    .A2(_1287_),
    .B1(_1296_),
    .Y(_1305_));
 sky130_fd_sc_hd__nand2_1 _3557_ (.A(net272),
    .B(net138),
    .Y(_1315_));
 sky130_fd_sc_hd__o211a_1 _3558_ (.A1(_1315_),
    .A2(_1221_),
    .B1(_1296_),
    .C1(_1277_),
    .X(_1326_));
 sky130_fd_sc_hd__nand2_1 _3559_ (.A(net312),
    .B(net132),
    .Y(_1336_));
 sky130_fd_sc_hd__nand4_2 _3560_ (.A(net119),
    .B(net336),
    .C(net323),
    .D(net125),
    .Y(_1347_));
 sky130_fd_sc_hd__a22oi_4 _3561_ (.A1(net119),
    .A2(net332),
    .B1(net324),
    .B2(net125),
    .Y(_1358_));
 sky130_fd_sc_hd__a21oi_2 _3562_ (.A1(_1336_),
    .A2(_1347_),
    .B1(_1358_),
    .Y(_1368_));
 sky130_fd_sc_hd__o21bai_4 _3563_ (.A1(_1305_),
    .A2(_1326_),
    .B1_N(_1368_),
    .Y(_1379_));
 sky130_fd_sc_hd__nand2_2 _3564_ (.A(net259),
    .B(net151),
    .Y(_1390_));
 sky130_fd_sc_hd__a21oi_1 _3565_ (.A1(_1277_),
    .A2(_1287_),
    .B1(_1390_),
    .Y(_1401_));
 sky130_fd_sc_hd__inv_4 _3566_ (.A(net259),
    .Y(_1412_));
 sky130_fd_sc_hd__clkbuf_8 _3567_ (.A(_1412_),
    .X(_1423_));
 sky130_fd_sc_hd__inv_2 _3568_ (.A(net154),
    .Y(_1434_));
 sky130_fd_sc_hd__buf_4 _3569_ (.A(_1434_),
    .X(_1445_));
 sky130_fd_sc_hd__o221a_1 _3570_ (.A1(_1423_),
    .A2(_1445_),
    .B1(_1315_),
    .B2(_1221_),
    .C1(_1277_),
    .X(_1456_));
 sky130_fd_sc_hd__o21ai_2 _3571_ (.A1(_1401_),
    .A2(_1456_),
    .B1(_1368_),
    .Y(_1466_));
 sky130_fd_sc_hd__a21boi_4 _3572_ (.A1(_1249_),
    .A2(_1379_),
    .B1_N(_1466_),
    .Y(_1477_));
 sky130_fd_sc_hd__a21o_1 _3573_ (.A1(_1165_),
    .A2(_1193_),
    .B1(_1477_),
    .X(_1488_));
 sky130_fd_sc_hd__and2_1 _3574_ (.A(net144),
    .B(net138),
    .X(_1499_));
 sky130_fd_sc_hd__a32o_1 _3575_ (.A1(net283),
    .A2(net272),
    .A3(_1499_),
    .B1(_1296_),
    .B2(_1277_),
    .X(_1510_));
 sky130_fd_sc_hd__nand2_1 _3576_ (.A(net259),
    .B(net145),
    .Y(_1521_));
 sky130_fd_sc_hd__nand2_1 _3577_ (.A(_1521_),
    .B(_1315_),
    .Y(_1531_));
 sky130_fd_sc_hd__nand4_1 _3578_ (.A(net272),
    .B(net260),
    .C(net145),
    .D(net138),
    .Y(_1542_));
 sky130_fd_sc_hd__a21oi_1 _3579_ (.A1(_1531_),
    .A2(_1542_),
    .B1(_1296_),
    .Y(_1553_));
 sky130_fd_sc_hd__and3_1 _3580_ (.A(_1531_),
    .B(_1542_),
    .C(_1296_),
    .X(_1564_));
 sky130_fd_sc_hd__nand2_1 _3581_ (.A(net312),
    .B(net125),
    .Y(_1575_));
 sky130_fd_sc_hd__nand2_1 _3582_ (.A(net119),
    .B(net321),
    .Y(_1586_));
 sky130_fd_sc_hd__nand4_4 _3583_ (.A(\mixer_q.nco_reg[8] ),
    .B(net321),
    .C(net312),
    .D(net125),
    .Y(_1597_));
 sky130_fd_sc_hd__nand2_1 _3584_ (.A(net296),
    .B(net131),
    .Y(_1607_));
 sky130_fd_sc_hd__a22oi_2 _3585_ (.A1(_1575_),
    .A2(_1586_),
    .B1(_1597_),
    .B2(_1607_),
    .Y(_1618_));
 sky130_fd_sc_hd__o21bai_2 _3586_ (.A1(_1553_),
    .A2(_1564_),
    .B1_N(_1618_),
    .Y(_1629_));
 sky130_fd_sc_hd__nand4_1 _3587_ (.A(_1531_),
    .B(_1542_),
    .C(net259),
    .D(net151),
    .Y(_1640_));
 sky130_fd_sc_hd__nand3b_2 _3588_ (.A_N(_1553_),
    .B(_1640_),
    .C(_1618_),
    .Y(_1651_));
 sky130_fd_sc_hd__a21bo_4 _3589_ (.A1(_1510_),
    .A2(_1629_),
    .B1_N(_1651_),
    .X(_1662_));
 sky130_fd_sc_hd__o311a_1 _3590_ (.A1(net170),
    .A2(net164),
    .A3(net157),
    .B1(_1662_),
    .C1(net258),
    .X(_1673_));
 sky130_fd_sc_hd__o31a_2 _3591_ (.A1(net170),
    .A2(net164),
    .A3(net157),
    .B1(net258),
    .X(_1684_));
 sky130_fd_sc_hd__nor2_1 _3592_ (.A(_1684_),
    .B(_1662_),
    .Y(_1695_));
 sky130_fd_sc_hd__nand3_4 _3593_ (.A(net101),
    .B(net106),
    .C(net346),
    .Y(_1705_));
 sky130_fd_sc_hd__nand2_1 _3594_ (.A(net112),
    .B(net333),
    .Y(_1716_));
 sky130_fd_sc_hd__clkinv_4 _3595_ (.A(net364),
    .Y(_1727_));
 sky130_fd_sc_hd__a22oi_4 _3596_ (.A1(net106),
    .A2(net346),
    .B1(_1727_),
    .B2(net101),
    .Y(_1738_));
 sky130_fd_sc_hd__o22ai_4 _3597_ (.A1(net358),
    .A2(_1705_),
    .B1(_1716_),
    .B2(_1738_),
    .Y(_1749_));
 sky130_fd_sc_hd__inv_2 _3598_ (.A(net111),
    .Y(_1760_));
 sky130_fd_sc_hd__buf_4 _3599_ (.A(_1760_),
    .X(_1771_));
 sky130_fd_sc_hd__inv_6 _3600_ (.A(net323),
    .Y(_1782_));
 sky130_fd_sc_hd__buf_6 _3601_ (.A(_1782_),
    .X(_1793_));
 sky130_fd_sc_hd__nand3_4 _3602_ (.A(net100),
    .B(net107),
    .C(net332),
    .Y(_1804_));
 sky130_fd_sc_hd__nor2_1 _3603_ (.A(net340),
    .B(_1804_),
    .Y(_1815_));
 sky130_fd_sc_hd__clkinv_4 _3604_ (.A(net347),
    .Y(_1825_));
 sky130_fd_sc_hd__a22oi_4 _3605_ (.A1(net107),
    .A2(net332),
    .B1(_1825_),
    .B2(net101),
    .Y(_1836_));
 sky130_fd_sc_hd__o22ai_4 _3606_ (.A1(_1771_),
    .A2(net96),
    .B1(_1815_),
    .B2(_1836_),
    .Y(_1847_));
 sky130_fd_sc_hd__clkinv_8 _3607_ (.A(net100),
    .Y(_1858_));
 sky130_fd_sc_hd__buf_6 _3608_ (.A(_1858_),
    .X(_1869_));
 sky130_fd_sc_hd__o2bb2ai_2 _3609_ (.A1_N(net107),
    .A2_N(net332),
    .B1(net346),
    .B2(_1869_),
    .Y(_1880_));
 sky130_fd_sc_hd__o2111ai_4 _3610_ (.A1(net346),
    .A2(_1804_),
    .B1(net321),
    .C1(net112),
    .D1(_1880_),
    .Y(_1891_));
 sky130_fd_sc_hd__nand3_2 _3611_ (.A(_1749_),
    .B(_1847_),
    .C(_1891_),
    .Y(_1902_));
 sky130_fd_sc_hd__nand2_1 _3612_ (.A(net115),
    .B(net321),
    .Y(_1913_));
 sky130_fd_sc_hd__o21bai_1 _3613_ (.A1(_1815_),
    .A2(_1836_),
    .B1_N(_1913_),
    .Y(_1924_));
 sky130_fd_sc_hd__o2bb2ai_4 _3614_ (.A1_N(net106),
    .A2_N(net346),
    .B1(net358),
    .B2(_1869_),
    .Y(_1934_));
 sky130_fd_sc_hd__and2_1 _3615_ (.A(net112),
    .B(net333),
    .X(_1945_));
 sky130_fd_sc_hd__nor2_1 _3616_ (.A(net358),
    .B(_1705_),
    .Y(_1956_));
 sky130_fd_sc_hd__a21oi_1 _3617_ (.A1(_1934_),
    .A2(_1945_),
    .B1(_1956_),
    .Y(_1967_));
 sky130_fd_sc_hd__o221ai_2 _3618_ (.A1(_1771_),
    .A2(net96),
    .B1(_1804_),
    .B2(net346),
    .C1(_1880_),
    .Y(_1978_));
 sky130_fd_sc_hd__nand3_2 _3619_ (.A(_1924_),
    .B(_1967_),
    .C(_1978_),
    .Y(_1989_));
 sky130_fd_sc_hd__nand4_2 _3620_ (.A(net296),
    .B(net117),
    .C(net312),
    .D(net123),
    .Y(_2000_));
 sky130_fd_sc_hd__nand2_1 _3621_ (.A(net119),
    .B(net312),
    .Y(_2011_));
 sky130_fd_sc_hd__nand2_1 _3622_ (.A(net296),
    .B(net128),
    .Y(_2022_));
 sky130_fd_sc_hd__nand2_1 _3623_ (.A(net283),
    .B(net131),
    .Y(_2033_));
 sky130_fd_sc_hd__a21oi_2 _3624_ (.A1(_2011_),
    .A2(_2022_),
    .B1(_2033_),
    .Y(_2044_));
 sky130_fd_sc_hd__nand2_1 _3625_ (.A(_2011_),
    .B(_2022_),
    .Y(_2054_));
 sky130_fd_sc_hd__a22oi_4 _3626_ (.A1(net283),
    .A2(net131),
    .B1(_2000_),
    .B2(_2054_),
    .Y(_2065_));
 sky130_fd_sc_hd__a21o_1 _3627_ (.A1(_2000_),
    .A2(_2044_),
    .B1(_2065_),
    .X(_2076_));
 sky130_fd_sc_hd__a21o_1 _3628_ (.A1(_1902_),
    .A2(_1989_),
    .B1(_2076_),
    .X(_2087_));
 sky130_fd_sc_hd__o21ai_2 _3629_ (.A1(_1956_),
    .A2(_1738_),
    .B1(_1945_),
    .Y(_2098_));
 sky130_fd_sc_hd__buf_6 _3630_ (.A(_1760_),
    .X(_2109_));
 sky130_fd_sc_hd__inv_4 _3631_ (.A(net337),
    .Y(_2120_));
 sky130_fd_sc_hd__o221ai_4 _3632_ (.A1(_2109_),
    .A2(_2120_),
    .B1(_1705_),
    .B2(net358),
    .C1(_1934_),
    .Y(_2131_));
 sky130_fd_sc_hd__o2bb2ai_4 _3633_ (.A1_N(net106),
    .A2_N(net358),
    .B1(net372),
    .B2(_1858_),
    .Y(_2142_));
 sky130_fd_sc_hd__nand3_4 _3634_ (.A(net101),
    .B(net106),
    .C(net358),
    .Y(_2153_));
 sky130_fd_sc_hd__nand2_1 _3635_ (.A(net112),
    .B(net346),
    .Y(_2163_));
 sky130_fd_sc_hd__o21ai_1 _3636_ (.A1(net372),
    .A2(_2153_),
    .B1(_2163_),
    .Y(_2174_));
 sky130_fd_sc_hd__nand2_1 _3637_ (.A(_2142_),
    .B(_2174_),
    .Y(_2185_));
 sky130_fd_sc_hd__nand3_4 _3638_ (.A(_2098_),
    .B(_2131_),
    .C(_2185_),
    .Y(_2196_));
 sky130_fd_sc_hd__o21ai_1 _3639_ (.A1(_1956_),
    .A2(_1738_),
    .B1(_1716_),
    .Y(_2207_));
 sky130_fd_sc_hd__inv_6 _3640_ (.A(net366),
    .Y(_2218_));
 sky130_fd_sc_hd__a22oi_4 _3641_ (.A1(net106),
    .A2(net358),
    .B1(_2218_),
    .B2(net101),
    .Y(_2229_));
 sky130_fd_sc_hd__o22ai_2 _3642_ (.A1(net372),
    .A2(_2153_),
    .B1(_2163_),
    .B2(_2229_),
    .Y(_2240_));
 sky130_fd_sc_hd__o2111ai_4 _3643_ (.A1(net358),
    .A2(_1705_),
    .B1(net332),
    .C1(net112),
    .D1(_1934_),
    .Y(_2251_));
 sky130_fd_sc_hd__nand3_4 _3644_ (.A(_2207_),
    .B(_2240_),
    .C(_2251_),
    .Y(_2261_));
 sky130_fd_sc_hd__nand2_1 _3645_ (.A(_1575_),
    .B(_1586_),
    .Y(_2272_));
 sky130_fd_sc_hd__a22o_1 _3646_ (.A1(net296),
    .A2(net131),
    .B1(_1597_),
    .B2(_2272_),
    .X(_2283_));
 sky130_fd_sc_hd__nand2_1 _3647_ (.A(net321),
    .B(net125),
    .Y(_2294_));
 sky130_fd_sc_hd__a21oi_1 _3648_ (.A1(_1575_),
    .A2(_1586_),
    .B1(_1607_),
    .Y(_2305_));
 sky130_fd_sc_hd__o21ai_1 _3649_ (.A1(_2011_),
    .A2(_2294_),
    .B1(_2305_),
    .Y(_2316_));
 sky130_fd_sc_hd__nand2_1 _3650_ (.A(_2283_),
    .B(_2316_),
    .Y(_2327_));
 sky130_fd_sc_hd__nand2_1 _3651_ (.A(_2261_),
    .B(_2327_),
    .Y(_2338_));
 sky130_fd_sc_hd__nand2_1 _3652_ (.A(_2196_),
    .B(_2338_),
    .Y(_2349_));
 sky130_fd_sc_hd__and4_1 _3653_ (.A(_2054_),
    .B(net131),
    .C(net283),
    .D(_2000_),
    .X(_2360_));
 sky130_fd_sc_hd__o211ai_2 _3654_ (.A1(_2360_),
    .A2(_2065_),
    .B1(_1989_),
    .C1(_1902_),
    .Y(_2370_));
 sky130_fd_sc_hd__and3_4 _3655_ (.A(_2087_),
    .B(_2349_),
    .C(_2370_),
    .X(_2381_));
 sky130_fd_sc_hd__a21oi_1 _3656_ (.A1(_1651_),
    .A2(_1629_),
    .B1(_1510_),
    .Y(_2392_));
 sky130_fd_sc_hd__nand3_2 _3657_ (.A(_1629_),
    .B(_1510_),
    .C(_1651_),
    .Y(_2403_));
 sky130_fd_sc_hd__inv_2 _3658_ (.A(_2403_),
    .Y(_2414_));
 sky130_fd_sc_hd__a22oi_4 _3659_ (.A1(net296),
    .A2(net131),
    .B1(_1597_),
    .B2(_2272_),
    .Y(_2425_));
 sky130_fd_sc_hd__a21oi_1 _3660_ (.A1(_1597_),
    .A2(_2305_),
    .B1(_2425_),
    .Y(_2436_));
 sky130_fd_sc_hd__nand2_1 _3661_ (.A(_2196_),
    .B(_2436_),
    .Y(_2447_));
 sky130_fd_sc_hd__nand2_1 _3662_ (.A(_2261_),
    .B(_2447_),
    .Y(_2458_));
 sky130_fd_sc_hd__a21oi_1 _3663_ (.A1(_2000_),
    .A2(_2044_),
    .B1(_2065_),
    .Y(_2468_));
 sky130_fd_sc_hd__nand3_1 _3664_ (.A(_1902_),
    .B(_1989_),
    .C(_2468_),
    .Y(_2479_));
 sky130_fd_sc_hd__o2bb2ai_1 _3665_ (.A1_N(_1902_),
    .A2_N(_1989_),
    .B1(_2065_),
    .B2(_2360_),
    .Y(_2490_));
 sky130_fd_sc_hd__nand3_4 _3666_ (.A(_2458_),
    .B(_2479_),
    .C(_2490_),
    .Y(_2501_));
 sky130_fd_sc_hd__o21a_2 _3667_ (.A1(_2392_),
    .A2(_2414_),
    .B1(_2501_),
    .X(_2512_));
 sky130_fd_sc_hd__and4_1 _3668_ (.A(net272),
    .B(net259),
    .C(net144),
    .D(net137),
    .X(_2523_));
 sky130_fd_sc_hd__and3_1 _3669_ (.A(_1531_),
    .B(net151),
    .C(net259),
    .X(_2534_));
 sky130_fd_sc_hd__and4_1 _3670_ (.A(net296),
    .B(net117),
    .C(net312),
    .D(net123),
    .X(_2545_));
 sky130_fd_sc_hd__nand2_4 _3671_ (.A(\mixer_q.nco_reg[4] ),
    .B(net143),
    .Y(_2555_));
 sky130_fd_sc_hd__o21a_1 _3672_ (.A1(net144),
    .A2(net137),
    .B1(net254),
    .X(_2566_));
 sky130_fd_sc_hd__o211ai_4 _3673_ (.A1(_1423_),
    .A2(_2555_),
    .B1(_2566_),
    .C1(net155),
    .Y(_2577_));
 sky130_fd_sc_hd__o21ai_2 _3674_ (.A1(net144),
    .A2(net137),
    .B1(net254),
    .Y(_2588_));
 sky130_fd_sc_hd__and3_1 _3675_ (.A(net253),
    .B(net144),
    .C(net137),
    .X(_2599_));
 sky130_fd_sc_hd__o21ai_4 _3676_ (.A1(_2588_),
    .A2(_2599_),
    .B1(_1390_),
    .Y(_2610_));
 sky130_fd_sc_hd__o211ai_4 _3677_ (.A1(_2545_),
    .A2(_2044_),
    .B1(_2577_),
    .C1(_2610_),
    .Y(_2621_));
 sky130_fd_sc_hd__nor2_1 _3678_ (.A(net144),
    .B(net137),
    .Y(_2631_));
 sky130_fd_sc_hd__nor3_2 _3679_ (.A(_1390_),
    .B(_2631_),
    .C(_1499_),
    .Y(_2642_));
 sky130_fd_sc_hd__buf_6 _3680_ (.A(_2642_),
    .X(_2653_));
 sky130_fd_sc_hd__nand3_2 _3681_ (.A(net254),
    .B(net144),
    .C(net137),
    .Y(_2664_));
 sky130_fd_sc_hd__a22oi_4 _3682_ (.A1(net254),
    .A2(net155),
    .B1(_2566_),
    .B2(_2664_),
    .Y(_2675_));
 sky130_fd_sc_hd__nor2_1 _3683_ (.A(_2545_),
    .B(_2044_),
    .Y(_2686_));
 sky130_fd_sc_hd__o21ai_4 _3684_ (.A1(_2653_),
    .A2(_2675_),
    .B1(_2686_),
    .Y(_2697_));
 sky130_fd_sc_hd__o211a_2 _3685_ (.A1(_2523_),
    .A2(_2534_),
    .B1(_2621_),
    .C1(_2697_),
    .X(_2707_));
 sky130_fd_sc_hd__a31o_2 _3686_ (.A1(net259),
    .A2(_1531_),
    .A3(net151),
    .B1(_2523_),
    .X(_2718_));
 sky130_fd_sc_hd__a21oi_4 _3687_ (.A1(_2621_),
    .A2(_2697_),
    .B1(_2718_),
    .Y(_2729_));
 sky130_fd_sc_hd__or2_1 _3688_ (.A(_2707_),
    .B(_2729_),
    .X(_2740_));
 sky130_fd_sc_hd__a21oi_4 _3689_ (.A1(_1847_),
    .A2(_1891_),
    .B1(_1749_),
    .Y(_2751_));
 sky130_fd_sc_hd__o21a_1 _3690_ (.A1(_2360_),
    .A2(_2065_),
    .B1(_1902_),
    .X(_2762_));
 sky130_fd_sc_hd__nand3_2 _3691_ (.A(net99),
    .B(net105),
    .C(net320),
    .Y(_2773_));
 sky130_fd_sc_hd__inv_6 _3692_ (.A(net307),
    .Y(_2783_));
 sky130_fd_sc_hd__buf_8 _3693_ (.A(_2783_),
    .X(_2794_));
 sky130_fd_sc_hd__nor2_1 _3694_ (.A(_2109_),
    .B(_2794_),
    .Y(_2805_));
 sky130_fd_sc_hd__o2bb2ai_4 _3695_ (.A1_N(net107),
    .A2_N(net321),
    .B1(net332),
    .B2(_1858_),
    .Y(_2816_));
 sky130_fd_sc_hd__o211a_1 _3696_ (.A1(net331),
    .A2(_2773_),
    .B1(_2805_),
    .C1(_2816_),
    .X(_2826_));
 sky130_fd_sc_hd__nand4_4 _3697_ (.A(_2120_),
    .B(net321),
    .C(net100),
    .D(net107),
    .Y(_2837_));
 sky130_fd_sc_hd__clkbuf_8 _3698_ (.A(_2783_),
    .X(_2848_));
 sky130_fd_sc_hd__o2bb2ai_4 _3699_ (.A1_N(_2816_),
    .A2_N(_2837_),
    .B1(_1771_),
    .B2(_2848_),
    .Y(_2859_));
 sky130_fd_sc_hd__o22ai_4 _3700_ (.A1(net341),
    .A2(_1804_),
    .B1(_1913_),
    .B2(_1836_),
    .Y(_2869_));
 sky130_fd_sc_hd__nand2_1 _3701_ (.A(_2859_),
    .B(_2869_),
    .Y(_2880_));
 sky130_fd_sc_hd__clkbuf_8 _3702_ (.A(_1782_),
    .X(_2886_));
 sky130_fd_sc_hd__o22a_1 _3703_ (.A1(net341),
    .A2(_1804_),
    .B1(_2886_),
    .B2(_1771_),
    .X(_2894_));
 sky130_fd_sc_hd__a21oi_1 _3704_ (.A1(_2816_),
    .A2(_2837_),
    .B1(_2805_),
    .Y(_2902_));
 sky130_fd_sc_hd__o22ai_4 _3705_ (.A1(_1836_),
    .A2(_2894_),
    .B1(_2826_),
    .B2(_2902_),
    .Y(_2909_));
 sky130_fd_sc_hd__a22oi_4 _3706_ (.A1(net295),
    .A2(net118),
    .B1(net124),
    .B2(net282),
    .Y(_2913_));
 sky130_fd_sc_hd__nand2_1 _3707_ (.A(net270),
    .B(net130),
    .Y(_2914_));
 sky130_fd_sc_hd__a41o_1 _3708_ (.A1(net295),
    .A2(net282),
    .A3(net117),
    .A4(net123),
    .B1(_2914_),
    .X(_2915_));
 sky130_fd_sc_hd__and4_1 _3709_ (.A(net295),
    .B(net282),
    .C(net117),
    .D(net123),
    .X(_2916_));
 sky130_fd_sc_hd__o21ai_2 _3710_ (.A1(_2913_),
    .A2(_2916_),
    .B1(_2914_),
    .Y(_2917_));
 sky130_fd_sc_hd__o21a_1 _3711_ (.A1(_2913_),
    .A2(_2915_),
    .B1(_2917_),
    .X(_2918_));
 sky130_fd_sc_hd__o211a_1 _3712_ (.A1(_2826_),
    .A2(_2880_),
    .B1(_2909_),
    .C1(_2918_),
    .X(_2919_));
 sky130_fd_sc_hd__buf_2 _3713_ (.A(_2109_),
    .X(_2920_));
 sky130_fd_sc_hd__nand3_2 _3714_ (.A(_2816_),
    .B(_2837_),
    .C(net312),
    .Y(_2921_));
 sky130_fd_sc_hd__o211ai_4 _3715_ (.A1(_2920_),
    .A2(_2921_),
    .B1(_2869_),
    .C1(_2859_),
    .Y(_2922_));
 sky130_fd_sc_hd__a21oi_4 _3716_ (.A1(_2922_),
    .A2(_2909_),
    .B1(_2918_),
    .Y(_2923_));
 sky130_fd_sc_hd__o22ai_4 _3717_ (.A1(_2751_),
    .A2(_2762_),
    .B1(_2919_),
    .B2(_2923_),
    .Y(_2924_));
 sky130_fd_sc_hd__a21oi_1 _3718_ (.A1(_1902_),
    .A2(_2076_),
    .B1(_2751_),
    .Y(_2925_));
 sky130_fd_sc_hd__o2111ai_4 _3719_ (.A1(_2915_),
    .A2(_2913_),
    .B1(_2917_),
    .C1(_2922_),
    .D1(_2909_),
    .Y(_2926_));
 sky130_fd_sc_hd__inv_6 _3720_ (.A(net271),
    .Y(_2927_));
 sky130_fd_sc_hd__buf_6 _3721_ (.A(_2927_),
    .X(_2928_));
 sky130_fd_sc_hd__buf_6 _3722_ (.A(_2928_),
    .X(_2929_));
 sky130_fd_sc_hd__inv_2 _3723_ (.A(net133),
    .Y(_2930_));
 sky130_fd_sc_hd__buf_4 _3724_ (.A(_2930_),
    .X(_2931_));
 sky130_fd_sc_hd__o22a_1 _3725_ (.A1(_2929_),
    .A2(_2931_),
    .B1(_2913_),
    .B2(_2916_),
    .X(_2932_));
 sky130_fd_sc_hd__nand4_1 _3726_ (.A(net295),
    .B(net282),
    .C(net118),
    .D(net124),
    .Y(_2933_));
 sky130_fd_sc_hd__and4b_1 _3727_ (.A_N(_2913_),
    .B(_2933_),
    .C(net270),
    .D(net130),
    .X(_2934_));
 sky130_fd_sc_hd__o211a_1 _3728_ (.A1(_2920_),
    .A2(_2921_),
    .B1(_2869_),
    .C1(_2859_),
    .X(_2935_));
 sky130_fd_sc_hd__o2111ai_2 _3729_ (.A1(net331),
    .A2(_2773_),
    .B1(net309),
    .C1(net111),
    .D1(_2816_),
    .Y(_2936_));
 sky130_fd_sc_hd__a2bb2oi_2 _3730_ (.A1_N(_1836_),
    .A2_N(_2894_),
    .B1(_2936_),
    .B2(_2859_),
    .Y(_2937_));
 sky130_fd_sc_hd__o22ai_4 _3731_ (.A1(_2932_),
    .A2(_2934_),
    .B1(_2935_),
    .B2(_2937_),
    .Y(_2938_));
 sky130_fd_sc_hd__nand3_2 _3732_ (.A(_2925_),
    .B(_2926_),
    .C(_2938_),
    .Y(_2939_));
 sky130_fd_sc_hd__nand3b_4 _3733_ (.A_N(_2740_),
    .B(_2924_),
    .C(_2939_),
    .Y(_2940_));
 sky130_fd_sc_hd__a2bb2oi_4 _3734_ (.A1_N(_2751_),
    .A2_N(_2762_),
    .B1(_2926_),
    .B2(_2938_),
    .Y(_2941_));
 sky130_fd_sc_hd__nand2_2 _3735_ (.A(_2925_),
    .B(_2926_),
    .Y(_2942_));
 sky130_fd_sc_hd__nor2_1 _3736_ (.A(_2923_),
    .B(_2942_),
    .Y(_2943_));
 sky130_fd_sc_hd__o22ai_4 _3737_ (.A1(_2707_),
    .A2(_2729_),
    .B1(_2941_),
    .B2(_2943_),
    .Y(_2944_));
 sky130_fd_sc_hd__a2bb2oi_4 _3738_ (.A1_N(_2381_),
    .A2_N(_2512_),
    .B1(_2940_),
    .B2(_2944_),
    .Y(_2945_));
 sky130_fd_sc_hd__inv_2 _3739_ (.A(_2501_),
    .Y(_2946_));
 sky130_fd_sc_hd__nand3_2 _3740_ (.A(_2087_),
    .B(_2349_),
    .C(_2370_),
    .Y(_2947_));
 sky130_fd_sc_hd__a21o_1 _3741_ (.A1(_1651_),
    .A2(_1629_),
    .B1(_1510_),
    .X(_2948_));
 sky130_fd_sc_hd__and3_1 _3742_ (.A(_2947_),
    .B(_2948_),
    .C(_2403_),
    .X(_2949_));
 sky130_fd_sc_hd__o211a_1 _3743_ (.A1(_2946_),
    .A2(_2949_),
    .B1(_2940_),
    .C1(_2944_),
    .X(_2950_));
 sky130_fd_sc_hd__o22ai_2 _3744_ (.A1(_1673_),
    .A2(_1695_),
    .B1(_2945_),
    .B2(_2950_),
    .Y(_2951_));
 sky130_fd_sc_hd__and3_1 _3745_ (.A(_1662_),
    .B(_1165_),
    .C(_1193_),
    .X(_2952_));
 sky130_fd_sc_hd__a21oi_2 _3746_ (.A1(_1165_),
    .A2(_1193_),
    .B1(_1662_),
    .Y(_2953_));
 sky130_fd_sc_hd__o221ai_4 _3747_ (.A1(_2923_),
    .A2(_2942_),
    .B1(_2729_),
    .B2(_2707_),
    .C1(_2924_),
    .Y(_2954_));
 sky130_fd_sc_hd__a21o_1 _3748_ (.A1(_2939_),
    .A2(_2924_),
    .B1(_2740_),
    .X(_2955_));
 sky130_fd_sc_hd__o211ai_4 _3749_ (.A1(_2381_),
    .A2(_2512_),
    .B1(_2954_),
    .C1(_2955_),
    .Y(_2956_));
 sky130_fd_sc_hd__o211ai_4 _3750_ (.A1(_2946_),
    .A2(_2949_),
    .B1(_2940_),
    .C1(_2944_),
    .Y(_2957_));
 sky130_fd_sc_hd__o211ai_2 _3751_ (.A1(_2952_),
    .A2(_2953_),
    .B1(_2956_),
    .C1(_2957_),
    .Y(_2958_));
 sky130_fd_sc_hd__nand3_1 _3752_ (.A(_2501_),
    .B(_2948_),
    .C(_2403_),
    .Y(_2959_));
 sky130_fd_sc_hd__a21o_1 _3753_ (.A1(_1466_),
    .A2(_1379_),
    .B1(_1249_),
    .X(_2960_));
 sky130_fd_sc_hd__nand3_1 _3754_ (.A(_1249_),
    .B(_1466_),
    .C(_1379_),
    .Y(_2961_));
 sky130_fd_sc_hd__nand2_1 _3755_ (.A(_2960_),
    .B(_2961_),
    .Y(_2962_));
 sky130_fd_sc_hd__and4b_1 _3756_ (.A_N(net371),
    .B(net359),
    .C(net101),
    .D(net106),
    .X(_2963_));
 sky130_fd_sc_hd__o21bai_4 _3757_ (.A1(_2229_),
    .A2(_2963_),
    .B1_N(_2163_),
    .Y(_2964_));
 sky130_fd_sc_hd__buf_6 _3758_ (.A(_1825_),
    .X(_2965_));
 sky130_fd_sc_hd__o221ai_4 _3759_ (.A1(_2109_),
    .A2(_2965_),
    .B1(_2153_),
    .B2(net371),
    .C1(_2142_),
    .Y(_2966_));
 sky130_fd_sc_hd__o2bb2ai_4 _3760_ (.A1_N(net106),
    .A2_N(net372),
    .B1(net382),
    .B2(_1858_),
    .Y(_2967_));
 sky130_fd_sc_hd__and2_2 _3761_ (.A(net113),
    .B(net362),
    .X(_2968_));
 sky130_fd_sc_hd__nand3_4 _3762_ (.A(net101),
    .B(net108),
    .C(net372),
    .Y(_2969_));
 sky130_fd_sc_hd__nor2_2 _3763_ (.A(net382),
    .B(_2969_),
    .Y(_2970_));
 sky130_fd_sc_hd__a21oi_4 _3764_ (.A1(_2967_),
    .A2(_2968_),
    .B1(_2970_),
    .Y(_2971_));
 sky130_fd_sc_hd__nand3_4 _3765_ (.A(_2964_),
    .B(_2966_),
    .C(_2971_),
    .Y(_2972_));
 sky130_fd_sc_hd__buf_6 _3766_ (.A(_2794_),
    .X(_2973_));
 sky130_fd_sc_hd__nand2_4 _3767_ (.A(net119),
    .B(net334),
    .Y(_2974_));
 sky130_fd_sc_hd__nor2_1 _3768_ (.A(_2294_),
    .B(_2974_),
    .Y(_2975_));
 sky130_fd_sc_hd__o22a_1 _3769_ (.A1(_2973_),
    .A2(_2931_),
    .B1(_1358_),
    .B2(_2975_),
    .X(_2976_));
 sky130_fd_sc_hd__a22o_1 _3770_ (.A1(net121),
    .A2(net336),
    .B1(net323),
    .B2(net127),
    .X(_2977_));
 sky130_fd_sc_hd__and4_2 _3771_ (.A(_2977_),
    .B(_1347_),
    .C(net311),
    .D(net132),
    .X(_2978_));
 sky130_fd_sc_hd__o21ai_1 _3772_ (.A1(_2229_),
    .A2(_2963_),
    .B1(_2163_),
    .Y(_2979_));
 sky130_fd_sc_hd__o2111ai_4 _3773_ (.A1(net371),
    .A2(_2153_),
    .B1(net346),
    .C1(net112),
    .D1(_2142_),
    .Y(_2980_));
 sky130_fd_sc_hd__nand2_2 _3774_ (.A(net113),
    .B(net361),
    .Y(_2981_));
 sky130_fd_sc_hd__inv_6 _3775_ (.A(net381),
    .Y(_2982_));
 sky130_fd_sc_hd__a22oi_4 _3776_ (.A1(net108),
    .A2(net371),
    .B1(_2982_),
    .B2(net101),
    .Y(_2983_));
 sky130_fd_sc_hd__o22ai_2 _3777_ (.A1(net382),
    .A2(_2969_),
    .B1(_2981_),
    .B2(_2983_),
    .Y(_2984_));
 sky130_fd_sc_hd__nand3_4 _3778_ (.A(_2979_),
    .B(_2980_),
    .C(_2984_),
    .Y(_2985_));
 sky130_fd_sc_hd__o21ai_1 _3779_ (.A1(_2976_),
    .A2(_2978_),
    .B1(_2985_),
    .Y(_2986_));
 sky130_fd_sc_hd__and4_1 _3780_ (.A(_2272_),
    .B(net131),
    .C(net296),
    .D(_1597_),
    .X(_2987_));
 sky130_fd_sc_hd__o2bb2ai_2 _3781_ (.A1_N(_2261_),
    .A2_N(_2196_),
    .B1(_2425_),
    .B2(_2987_),
    .Y(_2988_));
 sky130_fd_sc_hd__nand4_1 _3782_ (.A(_2261_),
    .B(_2196_),
    .C(_2283_),
    .D(_2316_),
    .Y(_2989_));
 sky130_fd_sc_hd__a22oi_2 _3783_ (.A1(_2972_),
    .A2(_2986_),
    .B1(_2988_),
    .B2(_2989_),
    .Y(_2990_));
 sky130_fd_sc_hd__a21oi_1 _3784_ (.A1(_2098_),
    .A2(_2131_),
    .B1(_2185_),
    .Y(_2991_));
 sky130_fd_sc_hd__a21oi_2 _3785_ (.A1(_2964_),
    .A2(_2966_),
    .B1(_2971_),
    .Y(_2992_));
 sky130_fd_sc_hd__o21ai_1 _3786_ (.A1(_1358_),
    .A2(_2975_),
    .B1(_1336_),
    .Y(_2993_));
 sky130_fd_sc_hd__nand4_1 _3787_ (.A(_2977_),
    .B(_1347_),
    .C(net311),
    .D(net132),
    .Y(_2994_));
 sky130_fd_sc_hd__nand2_1 _3788_ (.A(_2993_),
    .B(_2994_),
    .Y(_2995_));
 sky130_fd_sc_hd__a31oi_2 _3789_ (.A1(_2964_),
    .A2(_2966_),
    .A3(_2971_),
    .B1(_2995_),
    .Y(_2996_));
 sky130_fd_sc_hd__o221ai_4 _3790_ (.A1(_2991_),
    .A2(_2447_),
    .B1(_2992_),
    .B2(_2996_),
    .C1(_2988_),
    .Y(_2997_));
 sky130_fd_sc_hd__o21ai_1 _3791_ (.A1(_2962_),
    .A2(_2990_),
    .B1(_2997_),
    .Y(_2998_));
 sky130_fd_sc_hd__o2bb2ai_1 _3792_ (.A1_N(_2947_),
    .A2_N(_2501_),
    .B1(_2392_),
    .B2(_2414_),
    .Y(_2999_));
 sky130_fd_sc_hd__o211ai_2 _3793_ (.A1(_2381_),
    .A2(_2959_),
    .B1(_2998_),
    .C1(_2999_),
    .Y(_3000_));
 sky130_fd_sc_hd__o21a_1 _3794_ (.A1(_2962_),
    .A2(_2990_),
    .B1(_2997_),
    .X(_3001_));
 sky130_fd_sc_hd__o211ai_1 _3795_ (.A1(_2392_),
    .A2(_2414_),
    .B1(_2947_),
    .C1(_2501_),
    .Y(_3002_));
 sky130_fd_sc_hd__nand2_1 _3796_ (.A(_2948_),
    .B(_2403_),
    .Y(_3003_));
 sky130_fd_sc_hd__a21o_1 _3797_ (.A1(_2947_),
    .A2(_2501_),
    .B1(_3003_),
    .X(_3004_));
 sky130_fd_sc_hd__nand3_2 _3798_ (.A(_3001_),
    .B(_3002_),
    .C(_3004_),
    .Y(_3005_));
 sky130_fd_sc_hd__a21oi_2 _3799_ (.A1(_1156_),
    .A2(_1183_),
    .B1(_1477_),
    .Y(_3006_));
 sky130_fd_sc_hd__and3_1 _3800_ (.A(_1156_),
    .B(_1477_),
    .C(_1183_),
    .X(_3007_));
 sky130_fd_sc_hd__nor2_1 _3801_ (.A(_3006_),
    .B(_3007_),
    .Y(_3008_));
 sky130_fd_sc_hd__nand2_1 _3802_ (.A(_3005_),
    .B(_3008_),
    .Y(_3009_));
 sky130_fd_sc_hd__nand2_1 _3803_ (.A(_3000_),
    .B(_3009_),
    .Y(_3010_));
 sky130_fd_sc_hd__nand3_4 _3804_ (.A(_2951_),
    .B(_2958_),
    .C(_3010_),
    .Y(_3011_));
 sky130_fd_sc_hd__o22ai_1 _3805_ (.A1(_2952_),
    .A2(_2953_),
    .B1(_2945_),
    .B2(_2950_),
    .Y(_3012_));
 sky130_fd_sc_hd__o211a_1 _3806_ (.A1(_2381_),
    .A2(_2959_),
    .B1(_2998_),
    .C1(_2999_),
    .X(_3013_));
 sky130_fd_sc_hd__o21ai_1 _3807_ (.A1(_3013_),
    .A2(_3008_),
    .B1(_3005_),
    .Y(_3014_));
 sky130_fd_sc_hd__nand2_1 _3808_ (.A(_3012_),
    .B(_3014_),
    .Y(_3015_));
 sky130_fd_sc_hd__nor2_1 _3809_ (.A(_2952_),
    .B(_2953_),
    .Y(_3016_));
 sky130_fd_sc_hd__and3_1 _3810_ (.A(_2957_),
    .B(_3016_),
    .C(_2956_),
    .X(_3017_));
 sky130_fd_sc_hd__o2bb2ai_2 _3811_ (.A1_N(_1488_),
    .A2_N(_3011_),
    .B1(_3015_),
    .B2(_3017_),
    .Y(_3018_));
 sky130_fd_sc_hd__a21oi_2 _3812_ (.A1(_2957_),
    .A2(_3016_),
    .B1(_2945_),
    .Y(_3019_));
 sky130_fd_sc_hd__a21oi_2 _3813_ (.A1(_2939_),
    .A2(_2740_),
    .B1(_2941_),
    .Y(_3020_));
 sky130_fd_sc_hd__clkinv_4 _3814_ (.A(net304),
    .Y(_3021_));
 sky130_fd_sc_hd__clkbuf_8 _3815_ (.A(_3021_),
    .X(_3022_));
 sky130_fd_sc_hd__nand3_2 _3816_ (.A(net99),
    .B(net104),
    .C(net309),
    .Y(_3023_));
 sky130_fd_sc_hd__nor2_1 _3817_ (.A(net320),
    .B(_3023_),
    .Y(_3024_));
 sky130_fd_sc_hd__a22oi_4 _3818_ (.A1(net104),
    .A2(net309),
    .B1(_1782_),
    .B2(net99),
    .Y(_3025_));
 sky130_fd_sc_hd__o22ai_4 _3819_ (.A1(_3022_),
    .A2(_1771_),
    .B1(_3024_),
    .B2(_3025_),
    .Y(_3026_));
 sky130_fd_sc_hd__o2bb2ai_1 _3820_ (.A1_N(net104),
    .A2_N(net309),
    .B1(net320),
    .B2(_1869_),
    .Y(_3027_));
 sky130_fd_sc_hd__o2111ai_4 _3821_ (.A1(net320),
    .A2(_3023_),
    .B1(net295),
    .C1(net111),
    .D1(_3027_),
    .Y(_3028_));
 sky130_fd_sc_hd__o22a_1 _3822_ (.A1(net331),
    .A2(_2773_),
    .B1(_2848_),
    .B2(_2109_),
    .X(_3029_));
 sky130_fd_sc_hd__o2bb2a_1 _3823_ (.A1_N(net104),
    .A2_N(net320),
    .B1(net331),
    .B2(_1869_),
    .X(_3030_));
 sky130_fd_sc_hd__o2bb2ai_2 _3824_ (.A1_N(_3026_),
    .A2_N(_3028_),
    .B1(_3029_),
    .B2(_3030_),
    .Y(_3031_));
 sky130_fd_sc_hd__o2bb2ai_1 _3825_ (.A1_N(_2805_),
    .A2_N(_2816_),
    .B1(net331),
    .B2(_2773_),
    .Y(_3032_));
 sky130_fd_sc_hd__nand3_2 _3826_ (.A(_3032_),
    .B(_3028_),
    .C(_3026_),
    .Y(_3033_));
 sky130_fd_sc_hd__nand4_1 _3827_ (.A(net282),
    .B(net270),
    .C(net116),
    .D(net122),
    .Y(_3034_));
 sky130_fd_sc_hd__a22o_1 _3828_ (.A1(net282),
    .A2(net116),
    .B1(net122),
    .B2(net270),
    .X(_3035_));
 sky130_fd_sc_hd__a22o_1 _3829_ (.A1(net253),
    .A2(net129),
    .B1(_3034_),
    .B2(_3035_),
    .X(_3036_));
 sky130_fd_sc_hd__nand4_1 _3830_ (.A(_3035_),
    .B(net129),
    .C(net253),
    .D(_3034_),
    .Y(_3037_));
 sky130_fd_sc_hd__nand2_1 _3831_ (.A(_3036_),
    .B(_3037_),
    .Y(_3038_));
 sky130_fd_sc_hd__a21o_1 _3832_ (.A1(_3031_),
    .A2(_3033_),
    .B1(_3038_),
    .X(_3039_));
 sky130_fd_sc_hd__o21ai_1 _3833_ (.A1(_2913_),
    .A2(_2915_),
    .B1(_2917_),
    .Y(_3040_));
 sky130_fd_sc_hd__a21o_1 _3834_ (.A1(_3040_),
    .A2(_2922_),
    .B1(_2937_),
    .X(_3041_));
 sky130_fd_sc_hd__nand3_1 _3835_ (.A(_3031_),
    .B(_3033_),
    .C(_3038_),
    .Y(_3042_));
 sky130_fd_sc_hd__nand3_4 _3836_ (.A(_3039_),
    .B(_3041_),
    .C(_3042_),
    .Y(_3043_));
 sky130_fd_sc_hd__nand2_1 _3837_ (.A(_3031_),
    .B(_3033_),
    .Y(_3044_));
 sky130_fd_sc_hd__nand2_1 _3838_ (.A(_3044_),
    .B(_3038_),
    .Y(_3045_));
 sky130_fd_sc_hd__nand4_2 _3839_ (.A(_3031_),
    .B(_3033_),
    .C(_3036_),
    .D(_3037_),
    .Y(_3046_));
 sky130_fd_sc_hd__a21oi_1 _3840_ (.A1(_2922_),
    .A2(_3040_),
    .B1(_2937_),
    .Y(_3047_));
 sky130_fd_sc_hd__nand3_4 _3841_ (.A(_3045_),
    .B(_3046_),
    .C(_3047_),
    .Y(_3048_));
 sky130_fd_sc_hd__buf_6 _3842_ (.A(_1434_),
    .X(_3049_));
 sky130_fd_sc_hd__buf_6 _3843_ (.A(_3049_),
    .X(_3050_));
 sky130_fd_sc_hd__o21a_1 _3844_ (.A1(_1499_),
    .A2(_2631_),
    .B1(_3050_),
    .X(_3051_));
 sky130_fd_sc_hd__o31ai_1 _3845_ (.A1(_1390_),
    .A2(_2631_),
    .A3(_1499_),
    .B1(net260),
    .Y(_3052_));
 sky130_fd_sc_hd__o21a_1 _3846_ (.A1(_2914_),
    .A2(_2913_),
    .B1(_2933_),
    .X(_3053_));
 sky130_fd_sc_hd__o21ai_1 _3847_ (.A1(_2653_),
    .A2(_2675_),
    .B1(_3053_),
    .Y(_3054_));
 sky130_fd_sc_hd__o31ai_1 _3848_ (.A1(_3051_),
    .A2(_3052_),
    .A3(_3053_),
    .B1(_3054_),
    .Y(_3055_));
 sky130_fd_sc_hd__o21ai_1 _3849_ (.A1(_2599_),
    .A2(_2653_),
    .B1(_3055_),
    .Y(_3056_));
 sky130_fd_sc_hd__nor3_2 _3850_ (.A(_2642_),
    .B(_2675_),
    .C(_3053_),
    .Y(_3057_));
 sky130_fd_sc_hd__buf_8 _3851_ (.A(_1423_),
    .X(_3058_));
 sky130_fd_sc_hd__o22a_2 _3852_ (.A1(_3058_),
    .A2(_2555_),
    .B1(_2588_),
    .B2(_3050_),
    .X(_3059_));
 sky130_fd_sc_hd__nand3b_1 _3853_ (.A_N(_3057_),
    .B(_3054_),
    .C(_3059_),
    .Y(_3060_));
 sky130_fd_sc_hd__nand2_2 _3854_ (.A(_3056_),
    .B(_3060_),
    .Y(_3061_));
 sky130_fd_sc_hd__a21o_1 _3855_ (.A1(_3043_),
    .A2(_3048_),
    .B1(_3061_),
    .X(_3062_));
 sky130_fd_sc_hd__nand3_2 _3856_ (.A(_3043_),
    .B(_3048_),
    .C(_3061_),
    .Y(_3063_));
 sky130_fd_sc_hd__nand3_4 _3857_ (.A(_3020_),
    .B(_3062_),
    .C(_3063_),
    .Y(_3064_));
 sky130_fd_sc_hd__o22a_1 _3858_ (.A1(_2707_),
    .A2(_2729_),
    .B1(_2923_),
    .B2(_2942_),
    .X(_3065_));
 sky130_fd_sc_hd__a21oi_2 _3859_ (.A1(_3043_),
    .A2(_3048_),
    .B1(_3061_),
    .Y(_3066_));
 sky130_fd_sc_hd__and3_1 _3860_ (.A(_3043_),
    .B(_3048_),
    .C(_3061_),
    .X(_3067_));
 sky130_fd_sc_hd__o22ai_4 _3861_ (.A1(_2941_),
    .A2(_3065_),
    .B1(_3066_),
    .B2(_3067_),
    .Y(_3068_));
 sky130_fd_sc_hd__a21boi_4 _3862_ (.A1(_2697_),
    .A2(_2718_),
    .B1_N(_2621_),
    .Y(_3069_));
 sky130_fd_sc_hd__and3_1 _3863_ (.A(_3069_),
    .B(_1165_),
    .C(_1193_),
    .X(_3070_));
 sky130_fd_sc_hd__a21oi_4 _3864_ (.A1(_1165_),
    .A2(_1193_),
    .B1(_3069_),
    .Y(_3071_));
 sky130_fd_sc_hd__o2bb2ai_1 _3865_ (.A1_N(_3064_),
    .A2_N(_3068_),
    .B1(_3070_),
    .B2(_3071_),
    .Y(_3072_));
 sky130_fd_sc_hd__nor2_1 _3866_ (.A(_1684_),
    .B(_3069_),
    .Y(_3073_));
 sky130_fd_sc_hd__o311a_1 _3867_ (.A1(net170),
    .A2(net165),
    .A3(net158),
    .B1(_3069_),
    .C1(net258),
    .X(_3074_));
 sky130_fd_sc_hd__o211ai_2 _3868_ (.A1(_3073_),
    .A2(_3074_),
    .B1(_3064_),
    .C1(_3068_),
    .Y(_3075_));
 sky130_fd_sc_hd__nand3_4 _3869_ (.A(_3019_),
    .B(_3072_),
    .C(_3075_),
    .Y(_3076_));
 sky130_fd_sc_hd__o21ai_1 _3870_ (.A1(_3003_),
    .A2(_2381_),
    .B1(_2501_),
    .Y(_3077_));
 sky130_fd_sc_hd__nor2_1 _3871_ (.A(_1673_),
    .B(_1695_),
    .Y(_3078_));
 sky130_fd_sc_hd__a31oi_4 _3872_ (.A1(_2944_),
    .A2(_3077_),
    .A3(_2940_),
    .B1(_3078_),
    .Y(_3079_));
 sky130_fd_sc_hd__o211ai_4 _3873_ (.A1(_3071_),
    .A2(_3070_),
    .B1(_3068_),
    .C1(_3064_),
    .Y(_3080_));
 sky130_fd_sc_hd__o2bb2ai_2 _3874_ (.A1_N(_3064_),
    .A2_N(_3068_),
    .B1(_3073_),
    .B2(_3074_),
    .Y(_3081_));
 sky130_fd_sc_hd__o211ai_4 _3875_ (.A1(_2945_),
    .A2(_3079_),
    .B1(_3080_),
    .C1(_3081_),
    .Y(_3082_));
 sky130_fd_sc_hd__a22o_1 _3876_ (.A1(_1684_),
    .A2(_1662_),
    .B1(_3076_),
    .B2(_3082_),
    .X(_3083_));
 sky130_fd_sc_hd__o21a_4 _3877_ (.A1(net163),
    .A2(net157),
    .B1(net256),
    .X(_3084_));
 sky130_fd_sc_hd__and2_1 _3878_ (.A(net256),
    .B(net170),
    .X(_3085_));
 sky130_fd_sc_hd__buf_6 _3879_ (.A(_3085_),
    .X(_3086_));
 sky130_fd_sc_hd__o2111ai_4 _3880_ (.A1(_3084_),
    .A2(_3086_),
    .B1(_1662_),
    .C1(_3082_),
    .D1(_3076_),
    .Y(_3087_));
 sky130_fd_sc_hd__nand3b_4 _3881_ (.A_N(_3018_),
    .B(_3083_),
    .C(_3087_),
    .Y(_3088_));
 sky130_fd_sc_hd__inv_2 _3882_ (.A(_3088_),
    .Y(_3089_));
 sky130_fd_sc_hd__a21bo_1 _3883_ (.A1(_1202_),
    .A2(_1240_),
    .B1_N(_1212_),
    .X(_3090_));
 sky130_fd_sc_hd__nand4_1 _3884_ (.A(_1240_),
    .B(net152),
    .C(net273),
    .D(_1202_),
    .Y(_3091_));
 sky130_fd_sc_hd__nand2_2 _3885_ (.A(net348),
    .B(net127),
    .Y(_3092_));
 sky130_fd_sc_hd__clkbuf_4 _3886_ (.A(_3092_),
    .X(_3093_));
 sky130_fd_sc_hd__nand2_2 _3887_ (.A(net322),
    .B(net135),
    .Y(_3094_));
 sky130_fd_sc_hd__a22oi_4 _3888_ (.A1(net119),
    .A2(net348),
    .B1(net336),
    .B2(net125),
    .Y(_3095_));
 sky130_fd_sc_hd__o22ai_2 _3889_ (.A1(_2974_),
    .A2(_3093_),
    .B1(_3094_),
    .B2(_3095_),
    .Y(_3096_));
 sky130_fd_sc_hd__nand3_2 _3890_ (.A(_3090_),
    .B(_3091_),
    .C(_3096_),
    .Y(_3097_));
 sky130_fd_sc_hd__a21oi_1 _3891_ (.A1(_1202_),
    .A2(_1240_),
    .B1(_1212_),
    .Y(_3098_));
 sky130_fd_sc_hd__o211ai_2 _3892_ (.A1(_2928_),
    .A2(_3050_),
    .B1(_1202_),
    .C1(_1240_),
    .Y(_3099_));
 sky130_fd_sc_hd__o221ai_2 _3893_ (.A1(_3094_),
    .A2(_3095_),
    .B1(_3093_),
    .B2(_2974_),
    .C1(_3099_),
    .Y(_3100_));
 sky130_fd_sc_hd__nand2_1 _3894_ (.A(net297),
    .B(net146),
    .Y(_3101_));
 sky130_fd_sc_hd__nand2_1 _3895_ (.A(net310),
    .B(net140),
    .Y(_3102_));
 sky130_fd_sc_hd__nand2_2 _3896_ (.A(_3101_),
    .B(_3102_),
    .Y(_3103_));
 sky130_fd_sc_hd__and4_1 _3897_ (.A(net297),
    .B(net310),
    .C(net146),
    .D(net140),
    .X(_3104_));
 sky130_fd_sc_hd__a31o_1 _3898_ (.A1(net284),
    .A2(_3103_),
    .A3(net152),
    .B1(_3104_),
    .X(_3105_));
 sky130_fd_sc_hd__o211ai_1 _3899_ (.A1(_3098_),
    .A2(_3100_),
    .B1(_3105_),
    .C1(_3097_),
    .Y(_3106_));
 sky130_fd_sc_hd__o2bb2a_1 _3900_ (.A1_N(_3097_),
    .A2_N(_3106_),
    .B1(_3086_),
    .B2(_3084_),
    .X(_3107_));
 sky130_fd_sc_hd__o311a_1 _3901_ (.A1(net170),
    .A2(net164),
    .A3(net156),
    .B1(net258),
    .C1(_1477_),
    .X(_3108_));
 sky130_fd_sc_hd__nor2_1 _3902_ (.A(_1684_),
    .B(_1477_),
    .Y(_3109_));
 sky130_fd_sc_hd__o2bb2ai_1 _3903_ (.A1_N(_3000_),
    .A2_N(_3005_),
    .B1(_3108_),
    .B2(_3109_),
    .Y(_3110_));
 sky130_fd_sc_hd__nor2_1 _3904_ (.A(_2976_),
    .B(_2978_),
    .Y(_3111_));
 sky130_fd_sc_hd__a21oi_1 _3905_ (.A1(_3111_),
    .A2(_2972_),
    .B1(_2992_),
    .Y(_3112_));
 sky130_fd_sc_hd__a21o_1 _3906_ (.A1(_2261_),
    .A2(_2196_),
    .B1(_2327_),
    .X(_3113_));
 sky130_fd_sc_hd__o211ai_1 _3907_ (.A1(_2425_),
    .A2(_2987_),
    .B1(_2261_),
    .C1(_2196_),
    .Y(_3114_));
 sky130_fd_sc_hd__nand3_2 _3908_ (.A(_3112_),
    .B(_3113_),
    .C(_3114_),
    .Y(_3115_));
 sky130_fd_sc_hd__a21oi_1 _3909_ (.A1(_1466_),
    .A2(_1379_),
    .B1(_1249_),
    .Y(_3116_));
 sky130_fd_sc_hd__and3_1 _3910_ (.A(_1249_),
    .B(_1466_),
    .C(_1379_),
    .X(_3117_));
 sky130_fd_sc_hd__o2bb2ai_1 _3911_ (.A1_N(_3115_),
    .A2_N(_2997_),
    .B1(_3116_),
    .B2(_3117_),
    .Y(_3118_));
 sky130_fd_sc_hd__a21o_1 _3912_ (.A1(_1202_),
    .A2(_1240_),
    .B1(_1212_),
    .X(_3119_));
 sky130_fd_sc_hd__nand3b_1 _3913_ (.A_N(_3096_),
    .B(_3119_),
    .C(_3099_),
    .Y(_3120_));
 sky130_fd_sc_hd__a21oi_2 _3914_ (.A1(_3120_),
    .A2(_3097_),
    .B1(_3105_),
    .Y(_3121_));
 sky130_fd_sc_hd__o211a_1 _3915_ (.A1(_3098_),
    .A2(_3100_),
    .B1(_3105_),
    .C1(_3097_),
    .X(_3122_));
 sky130_fd_sc_hd__nor2_1 _3916_ (.A(_3121_),
    .B(_3122_),
    .Y(_3123_));
 sky130_fd_sc_hd__inv_4 _3917_ (.A(net396),
    .Y(_3124_));
 sky130_fd_sc_hd__clkbuf_8 _3918_ (.A(_3124_),
    .X(_3125_));
 sky130_fd_sc_hd__a21oi_2 _3919_ (.A1(net108),
    .A2(net382),
    .B1(_3125_),
    .Y(_3126_));
 sky130_fd_sc_hd__buf_4 _3920_ (.A(_1858_),
    .X(_3127_));
 sky130_fd_sc_hd__o221ai_4 _3921_ (.A1(_2109_),
    .A2(_1727_),
    .B1(_2969_),
    .B2(net382),
    .C1(_2967_),
    .Y(_3128_));
 sky130_fd_sc_hd__o21ai_4 _3922_ (.A1(_2983_),
    .A2(_2970_),
    .B1(_2968_),
    .Y(_3129_));
 sky130_fd_sc_hd__o211a_1 _3923_ (.A1(_3126_),
    .A2(_3127_),
    .B1(_3128_),
    .C1(_3129_),
    .X(_3130_));
 sky130_fd_sc_hd__nand2_1 _3924_ (.A(net108),
    .B(net383),
    .Y(_3131_));
 sky130_fd_sc_hd__a21oi_2 _3925_ (.A1(_3131_),
    .A2(net397),
    .B1(_3127_),
    .Y(_3132_));
 sky130_fd_sc_hd__o2111ai_4 _3926_ (.A1(net382),
    .A2(_2969_),
    .B1(net362),
    .C1(net113),
    .D1(_2967_),
    .Y(_3133_));
 sky130_fd_sc_hd__buf_8 _3927_ (.A(_1727_),
    .X(_3134_));
 sky130_fd_sc_hd__o22ai_4 _3928_ (.A1(_2109_),
    .A2(_3134_),
    .B1(_2983_),
    .B2(_2970_),
    .Y(_3135_));
 sky130_fd_sc_hd__a22o_1 _3929_ (.A1(net119),
    .A2(net348),
    .B1(net334),
    .B2(net125),
    .X(_3136_));
 sky130_fd_sc_hd__o221ai_4 _3930_ (.A1(_2886_),
    .A2(_2931_),
    .B1(_2974_),
    .B2(_3092_),
    .C1(_3136_),
    .Y(_3137_));
 sky130_fd_sc_hd__nor2_1 _3931_ (.A(_2974_),
    .B(_3092_),
    .Y(_3138_));
 sky130_fd_sc_hd__o21bai_2 _3932_ (.A1(_3095_),
    .A2(_3138_),
    .B1_N(_3094_),
    .Y(_3139_));
 sky130_fd_sc_hd__nand2_2 _3933_ (.A(_3137_),
    .B(_3139_),
    .Y(_3140_));
 sky130_fd_sc_hd__a31oi_2 _3934_ (.A1(_3132_),
    .A2(_3133_),
    .A3(_3135_),
    .B1(_3140_),
    .Y(_3141_));
 sky130_fd_sc_hd__o211ai_2 _3935_ (.A1(_2976_),
    .A2(_2978_),
    .B1(_2972_),
    .C1(_2985_),
    .Y(_3142_));
 sky130_fd_sc_hd__and3_1 _3936_ (.A(_1336_),
    .B(_2977_),
    .C(_1347_),
    .X(_3143_));
 sky130_fd_sc_hd__o211a_1 _3937_ (.A1(_1358_),
    .A2(_2975_),
    .B1(net311),
    .C1(net132),
    .X(_3144_));
 sky130_fd_sc_hd__o2bb2ai_1 _3938_ (.A1_N(_2972_),
    .A2_N(_2985_),
    .B1(_3143_),
    .B2(_3144_),
    .Y(_3145_));
 sky130_fd_sc_hd__o211ai_4 _3939_ (.A1(_3130_),
    .A2(_3141_),
    .B1(_3142_),
    .C1(_3145_),
    .Y(_3146_));
 sky130_fd_sc_hd__o211ai_4 _3940_ (.A1(_3143_),
    .A2(_3144_),
    .B1(_2972_),
    .C1(_2985_),
    .Y(_3147_));
 sky130_fd_sc_hd__inv_2 _3941_ (.A(_3147_),
    .Y(_3148_));
 sky130_fd_sc_hd__and3_2 _3942_ (.A(_3135_),
    .B(_3132_),
    .C(_3133_),
    .X(_3149_));
 sky130_fd_sc_hd__a21o_1 _3943_ (.A1(_3131_),
    .A2(net397),
    .B1(_3127_),
    .X(_3150_));
 sky130_fd_sc_hd__o21ai_1 _3944_ (.A1(_3095_),
    .A2(_3138_),
    .B1(_3094_),
    .Y(_3151_));
 sky130_fd_sc_hd__o2111ai_1 _3945_ (.A1(_2974_),
    .A2(_3093_),
    .B1(net322),
    .C1(net131),
    .D1(_3136_),
    .Y(_3152_));
 sky130_fd_sc_hd__nand2_1 _3946_ (.A(_3151_),
    .B(_3152_),
    .Y(_3153_));
 sky130_fd_sc_hd__a31oi_4 _3947_ (.A1(_3150_),
    .A2(_3129_),
    .A3(_3128_),
    .B1(_3153_),
    .Y(_3154_));
 sky130_fd_sc_hd__o2bb2ai_2 _3948_ (.A1_N(_2972_),
    .A2_N(_2985_),
    .B1(_2976_),
    .B2(_2978_),
    .Y(_3155_));
 sky130_fd_sc_hd__o21ai_4 _3949_ (.A1(_3149_),
    .A2(_3154_),
    .B1(_3155_),
    .Y(_3156_));
 sky130_fd_sc_hd__o2bb2ai_1 _3950_ (.A1_N(_3123_),
    .A2_N(_3146_),
    .B1(_3148_),
    .B2(_3156_),
    .Y(_3157_));
 sky130_fd_sc_hd__nand4_1 _3951_ (.A(_3115_),
    .B(_2997_),
    .C(_2960_),
    .D(_2961_),
    .Y(_3158_));
 sky130_fd_sc_hd__nand3_2 _3952_ (.A(_3118_),
    .B(_3157_),
    .C(_3158_),
    .Y(_3159_));
 sky130_fd_sc_hd__and3_1 _3953_ (.A(_1156_),
    .B(_3106_),
    .C(_1183_),
    .X(_3160_));
 sky130_fd_sc_hd__a21o_1 _3954_ (.A1(_3160_),
    .A2(_3097_),
    .B1(_3107_),
    .X(_3161_));
 sky130_fd_sc_hd__nand2_1 _3955_ (.A(_3146_),
    .B(_3123_),
    .Y(_3162_));
 sky130_fd_sc_hd__nand3_1 _3956_ (.A(_3115_),
    .B(_2997_),
    .C(_2962_),
    .Y(_3163_));
 sky130_fd_sc_hd__o211ai_4 _3957_ (.A1(_3148_),
    .A2(_3156_),
    .B1(_3162_),
    .C1(_3163_),
    .Y(_3164_));
 sky130_fd_sc_hd__a21oi_2 _3958_ (.A1(_3115_),
    .A2(_2997_),
    .B1(_2962_),
    .Y(_3165_));
 sky130_fd_sc_hd__o2bb2ai_1 _3959_ (.A1_N(_3159_),
    .A2_N(_3161_),
    .B1(_3164_),
    .B2(_3165_),
    .Y(_3166_));
 sky130_fd_sc_hd__o211ai_1 _3960_ (.A1(_3006_),
    .A2(_3007_),
    .B1(_3000_),
    .C1(_3005_),
    .Y(_3167_));
 sky130_fd_sc_hd__nand3_1 _3961_ (.A(_3110_),
    .B(_3166_),
    .C(_3167_),
    .Y(_3168_));
 sky130_fd_sc_hd__a2bb2oi_1 _3962_ (.A1_N(_3165_),
    .A2_N(_3164_),
    .B1(_3161_),
    .B2(_3159_),
    .Y(_3169_));
 sky130_fd_sc_hd__o2bb2ai_1 _3963_ (.A1_N(_3000_),
    .A2_N(_3005_),
    .B1(_3006_),
    .B2(_3007_),
    .Y(_3170_));
 sky130_fd_sc_hd__o211ai_2 _3964_ (.A1(_3013_),
    .A2(_3009_),
    .B1(_3169_),
    .C1(_3170_),
    .Y(_3171_));
 sky130_fd_sc_hd__a21boi_1 _3965_ (.A1(_3107_),
    .A2(_3168_),
    .B1_N(_3171_),
    .Y(_3172_));
 sky130_fd_sc_hd__o211ai_2 _3966_ (.A1(_3017_),
    .A2(_3015_),
    .B1(_3011_),
    .C1(_3006_),
    .Y(_3173_));
 sky130_fd_sc_hd__o211ai_1 _3967_ (.A1(_1673_),
    .A2(_1695_),
    .B1(_2956_),
    .C1(_2957_),
    .Y(_3174_));
 sky130_fd_sc_hd__nand3_1 _3968_ (.A(_3012_),
    .B(_3174_),
    .C(_3014_),
    .Y(_3175_));
 sky130_fd_sc_hd__clkbuf_8 _3969_ (.A(_3058_),
    .X(_3176_));
 sky130_fd_sc_hd__inv_4 _3970_ (.A(net173),
    .Y(_3177_));
 sky130_fd_sc_hd__buf_4 _3971_ (.A(_3177_),
    .X(_3178_));
 sky130_fd_sc_hd__o21a_2 _3972_ (.A1(_3176_),
    .A2(_3178_),
    .B1(_1183_),
    .X(_3179_));
 sky130_fd_sc_hd__o2bb2ai_1 _3973_ (.A1_N(_3011_),
    .A2_N(_3175_),
    .B1(_3179_),
    .B2(_1477_),
    .Y(_3180_));
 sky130_fd_sc_hd__nand3b_4 _3974_ (.A_N(_3172_),
    .B(_3173_),
    .C(_3180_),
    .Y(_3181_));
 sky130_fd_sc_hd__nand2_2 _3975_ (.A(net120),
    .B(net373),
    .Y(_3182_));
 sky130_fd_sc_hd__nand2_1 _3976_ (.A(net360),
    .B(net126),
    .Y(_3183_));
 sky130_fd_sc_hd__nand2_1 _3977_ (.A(_3182_),
    .B(_3183_),
    .Y(_3184_));
 sky130_fd_sc_hd__nand4_4 _3978_ (.A(net120),
    .B(net373),
    .C(net360),
    .D(net128),
    .Y(_3185_));
 sky130_fd_sc_hd__a22o_1 _3979_ (.A1(net349),
    .A2(net133),
    .B1(_3184_),
    .B2(_3185_),
    .X(_3186_));
 sky130_fd_sc_hd__nand4_2 _3980_ (.A(_3184_),
    .B(_3185_),
    .C(net349),
    .D(net133),
    .Y(_3187_));
 sky130_fd_sc_hd__and4_1 _3981_ (.A(net108),
    .B(net114),
    .C(net395),
    .D(net383),
    .X(_3188_));
 sky130_fd_sc_hd__a22oi_4 _3982_ (.A1(net108),
    .A2(net393),
    .B1(net384),
    .B2(net114),
    .Y(_3189_));
 sky130_fd_sc_hd__nor2_1 _3983_ (.A(_3188_),
    .B(_3189_),
    .Y(_3190_));
 sky130_fd_sc_hd__nand3_4 _3984_ (.A(_3186_),
    .B(_3187_),
    .C(_3190_),
    .Y(_3191_));
 sky130_fd_sc_hd__a22oi_4 _3985_ (.A1(net120),
    .A2(net374),
    .B1(net360),
    .B2(net126),
    .Y(_3192_));
 sky130_fd_sc_hd__nand2_2 _3986_ (.A(net349),
    .B(net133),
    .Y(_3193_));
 sky130_fd_sc_hd__o21ai_2 _3987_ (.A1(_3182_),
    .A2(_3183_),
    .B1(_3193_),
    .Y(_3194_));
 sky130_fd_sc_hd__a21o_1 _3988_ (.A1(_3184_),
    .A2(_3185_),
    .B1(_3193_),
    .X(_3195_));
 sky130_fd_sc_hd__o221ai_4 _3989_ (.A1(_3188_),
    .A2(_3189_),
    .B1(_3192_),
    .B2(_3194_),
    .C1(_3195_),
    .Y(_3196_));
 sky130_fd_sc_hd__nand4_4 _3990_ (.A(net121),
    .B(net383),
    .C(net373),
    .D(net126),
    .Y(_3197_));
 sky130_fd_sc_hd__nand2_1 _3991_ (.A(net373),
    .B(net127),
    .Y(_3198_));
 sky130_fd_sc_hd__nand2_1 _3992_ (.A(net121),
    .B(net384),
    .Y(_3199_));
 sky130_fd_sc_hd__nand2_1 _3993_ (.A(_3198_),
    .B(_3199_),
    .Y(_3200_));
 sky130_fd_sc_hd__o2bb2ai_2 _3994_ (.A1_N(_3197_),
    .A2_N(_3200_),
    .B1(_3134_),
    .B2(_2930_),
    .Y(_3201_));
 sky130_fd_sc_hd__nand4_2 _3995_ (.A(_3200_),
    .B(net133),
    .C(net360),
    .D(_3197_),
    .Y(_3202_));
 sky130_fd_sc_hd__nand2_1 _3996_ (.A(_3201_),
    .B(_3202_),
    .Y(_3203_));
 sky130_fd_sc_hd__nand2_4 _3997_ (.A(net114),
    .B(net393),
    .Y(_3204_));
 sky130_fd_sc_hd__o2bb2ai_4 _3998_ (.A1_N(_3191_),
    .A2_N(_3196_),
    .B1(_3203_),
    .B2(_3204_),
    .Y(_3205_));
 sky130_fd_sc_hd__nand4_4 _3999_ (.A(net336),
    .B(net323),
    .C(net146),
    .D(net140),
    .Y(_3206_));
 sky130_fd_sc_hd__nand2_1 _4000_ (.A(net335),
    .B(net139),
    .Y(_3207_));
 sky130_fd_sc_hd__nand2_1 _4001_ (.A(net323),
    .B(net146),
    .Y(_3208_));
 sky130_fd_sc_hd__nand2_2 _4002_ (.A(_3207_),
    .B(_3208_),
    .Y(_3209_));
 sky130_fd_sc_hd__o2bb2ai_1 _4003_ (.A1_N(_3206_),
    .A2_N(_3209_),
    .B1(_2848_),
    .B2(_1445_),
    .Y(_3210_));
 sky130_fd_sc_hd__nand2_1 _4004_ (.A(net360),
    .B(net133),
    .Y(_3211_));
 sky130_fd_sc_hd__a22oi_1 _4005_ (.A1(net120),
    .A2(net383),
    .B1(net373),
    .B2(net126),
    .Y(_3212_));
 sky130_fd_sc_hd__o21ai_1 _4006_ (.A1(_3211_),
    .A2(_3212_),
    .B1(_3197_),
    .Y(_3213_));
 sky130_fd_sc_hd__nand4_1 _4007_ (.A(_3209_),
    .B(net153),
    .C(net310),
    .D(_3206_),
    .Y(_3214_));
 sky130_fd_sc_hd__nand3_2 _4008_ (.A(_3210_),
    .B(_3213_),
    .C(_3214_),
    .Y(_3215_));
 sky130_fd_sc_hd__o21a_1 _4009_ (.A1(_3211_),
    .A2(_3212_),
    .B1(_3197_),
    .X(_3216_));
 sky130_fd_sc_hd__nand2_1 _4010_ (.A(net310),
    .B(net152),
    .Y(_3217_));
 sky130_fd_sc_hd__a21o_1 _4011_ (.A1(_3206_),
    .A2(_3209_),
    .B1(_3217_),
    .X(_3218_));
 sky130_fd_sc_hd__o211ai_4 _4012_ (.A1(_2794_),
    .A2(_3049_),
    .B1(_3206_),
    .C1(_3209_),
    .Y(_3219_));
 sky130_fd_sc_hd__nand3_1 _4013_ (.A(_3216_),
    .B(_3218_),
    .C(_3219_),
    .Y(_3220_));
 sky130_fd_sc_hd__buf_6 _4014_ (.A(_3220_),
    .X(_3221_));
 sky130_fd_sc_hd__nand2_1 _4015_ (.A(net323),
    .B(net153),
    .Y(_3222_));
 sky130_fd_sc_hd__nand4_4 _4016_ (.A(net349),
    .B(net335),
    .C(net147),
    .D(net140),
    .Y(_3223_));
 sky130_fd_sc_hd__a22oi_2 _4017_ (.A1(net335),
    .A2(net147),
    .B1(net139),
    .B2(net349),
    .Y(_3224_));
 sky130_fd_sc_hd__a21oi_2 _4018_ (.A1(_3222_),
    .A2(_3223_),
    .B1(_3224_),
    .Y(_3225_));
 sky130_fd_sc_hd__a21oi_1 _4019_ (.A1(_3215_),
    .A2(_3221_),
    .B1(_3225_),
    .Y(_3226_));
 sky130_fd_sc_hd__and3_1 _4020_ (.A(_3225_),
    .B(_3215_),
    .C(_3221_),
    .X(_3227_));
 sky130_fd_sc_hd__and2_2 _4021_ (.A(net113),
    .B(net393),
    .X(_3228_));
 sky130_fd_sc_hd__and3_1 _4022_ (.A(_3201_),
    .B(_3202_),
    .C(_3228_),
    .X(_3229_));
 sky130_fd_sc_hd__nand3_4 _4023_ (.A(_3229_),
    .B(_3196_),
    .C(_3191_),
    .Y(_3230_));
 sky130_fd_sc_hd__o21ai_2 _4024_ (.A1(_3226_),
    .A2(_3227_),
    .B1(_3230_),
    .Y(_3231_));
 sky130_fd_sc_hd__nand2_1 _4025_ (.A(net322),
    .B(net139),
    .Y(_3232_));
 sky130_fd_sc_hd__nand2_1 _4026_ (.A(net335),
    .B(net135),
    .Y(_3233_));
 sky130_fd_sc_hd__nand2_1 _4027_ (.A(_3232_),
    .B(_3233_),
    .Y(_3234_));
 sky130_fd_sc_hd__nand4_2 _4028_ (.A(net335),
    .B(net322),
    .C(net135),
    .D(net139),
    .Y(_3235_));
 sky130_fd_sc_hd__nand2_1 _4029_ (.A(net310),
    .B(net147),
    .Y(_3236_));
 sky130_fd_sc_hd__buf_4 _4030_ (.A(_3236_),
    .X(_3237_));
 sky130_fd_sc_hd__a21o_1 _4031_ (.A1(_3234_),
    .A2(_3235_),
    .B1(_3237_),
    .X(_3238_));
 sky130_fd_sc_hd__a21o_1 _4032_ (.A1(_3193_),
    .A2(_3185_),
    .B1(_3192_),
    .X(_3239_));
 sky130_fd_sc_hd__o211ai_2 _4033_ (.A1(_3094_),
    .A2(_3207_),
    .B1(_3234_),
    .C1(_3237_),
    .Y(_3240_));
 sky130_fd_sc_hd__a22oi_4 _4034_ (.A1(net322),
    .A2(net147),
    .B1(net139),
    .B2(net335),
    .Y(_3241_));
 sky130_fd_sc_hd__a21o_1 _4035_ (.A1(_3206_),
    .A2(_3217_),
    .B1(_3241_),
    .X(_3242_));
 sky130_fd_sc_hd__a31o_2 _4036_ (.A1(_3238_),
    .A2(_3239_),
    .A3(_3240_),
    .B1(_3242_),
    .X(_3243_));
 sky130_fd_sc_hd__a41o_1 _4037_ (.A1(net335),
    .A2(net322),
    .A3(net133),
    .A4(net139),
    .B1(_3236_),
    .X(_3244_));
 sky130_fd_sc_hd__a22oi_4 _4038_ (.A1(net335),
    .A2(net133),
    .B1(net139),
    .B2(net322),
    .Y(_3245_));
 sky130_fd_sc_hd__a21oi_2 _4039_ (.A1(_3193_),
    .A2(_3185_),
    .B1(_3192_),
    .Y(_3246_));
 sky130_fd_sc_hd__a21bo_1 _4040_ (.A1(_3234_),
    .A2(_3235_),
    .B1_N(_3237_),
    .X(_3247_));
 sky130_fd_sc_hd__o211a_1 _4041_ (.A1(_3244_),
    .A2(_3245_),
    .B1(_3246_),
    .C1(_3247_),
    .X(_3248_));
 sky130_fd_sc_hd__a21o_1 _4042_ (.A1(net102),
    .A2(net393),
    .B1(_3131_),
    .X(_3249_));
 sky130_fd_sc_hd__o211ai_1 _4043_ (.A1(net113),
    .A2(_3131_),
    .B1(net393),
    .C1(net102),
    .Y(_3250_));
 sky130_fd_sc_hd__o21ai_2 _4044_ (.A1(_3228_),
    .A2(_3249_),
    .B1(_3250_),
    .Y(_3251_));
 sky130_fd_sc_hd__a22oi_4 _4045_ (.A1(net113),
    .A2(net373),
    .B1(net360),
    .B2(net121),
    .Y(_3252_));
 sky130_fd_sc_hd__nor2_1 _4046_ (.A(_2981_),
    .B(_3182_),
    .Y(_3253_));
 sky130_fd_sc_hd__o21ai_4 _4047_ (.A1(_3252_),
    .A2(_3253_),
    .B1(_3093_),
    .Y(_3254_));
 sky130_fd_sc_hd__a22o_1 _4048_ (.A1(net113),
    .A2(net373),
    .B1(net360),
    .B2(net121),
    .X(_3255_));
 sky130_fd_sc_hd__nand4_4 _4049_ (.A(net114),
    .B(net121),
    .C(net373),
    .D(net360),
    .Y(_3256_));
 sky130_fd_sc_hd__nand4_4 _4050_ (.A(_3255_),
    .B(_3256_),
    .C(net349),
    .D(net127),
    .Y(_3257_));
 sky130_fd_sc_hd__nand3_4 _4051_ (.A(_3251_),
    .B(_3254_),
    .C(_3257_),
    .Y(_3258_));
 sky130_fd_sc_hd__nand4_1 _4052_ (.A(net102),
    .B(net109),
    .C(net393),
    .D(net383),
    .Y(_3259_));
 sky130_fd_sc_hd__a21oi_1 _4053_ (.A1(net113),
    .A2(net393),
    .B1(_3259_),
    .Y(_3260_));
 sky130_fd_sc_hd__a32oi_4 _4054_ (.A1(_3204_),
    .A2(net383),
    .A3(net108),
    .B1(net102),
    .B2(net393),
    .Y(_3261_));
 sky130_fd_sc_hd__o211ai_2 _4055_ (.A1(_2981_),
    .A2(_3182_),
    .B1(_3255_),
    .C1(_3093_),
    .Y(_3262_));
 sky130_fd_sc_hd__a21o_1 _4056_ (.A1(_3255_),
    .A2(_3256_),
    .B1(_3093_),
    .X(_3263_));
 sky130_fd_sc_hd__o211ai_4 _4057_ (.A1(_3260_),
    .A2(_3261_),
    .B1(_3262_),
    .C1(_3263_),
    .Y(_3264_));
 sky130_fd_sc_hd__o21a_1 _4058_ (.A1(_3192_),
    .A2(_3194_),
    .B1(_3195_),
    .X(_3265_));
 sky130_fd_sc_hd__a31o_1 _4059_ (.A1(net109),
    .A2(net383),
    .A3(_3228_),
    .B1(_3189_),
    .X(_3266_));
 sky130_fd_sc_hd__o2bb2ai_4 _4060_ (.A1_N(_3258_),
    .A2_N(_3264_),
    .B1(_3265_),
    .B2(_3266_),
    .Y(_3267_));
 sky130_fd_sc_hd__nand3b_4 _4061_ (.A_N(_3191_),
    .B(_3264_),
    .C(_3258_),
    .Y(_3268_));
 sky130_fd_sc_hd__nand3_1 _4062_ (.A(_3238_),
    .B(_3239_),
    .C(_3240_),
    .Y(_3269_));
 sky130_fd_sc_hd__clkbuf_4 _4063_ (.A(_3269_),
    .X(_3270_));
 sky130_fd_sc_hd__o211ai_4 _4064_ (.A1(_3244_),
    .A2(_3245_),
    .B1(_3246_),
    .C1(_3247_),
    .Y(_3271_));
 sky130_fd_sc_hd__buf_6 _4065_ (.A(_3271_),
    .X(_3272_));
 sky130_fd_sc_hd__a21oi_1 _4066_ (.A1(_3206_),
    .A2(_3217_),
    .B1(_3241_),
    .Y(_3273_));
 sky130_fd_sc_hd__a21o_1 _4067_ (.A1(_3270_),
    .A2(_3272_),
    .B1(_3273_),
    .X(_3274_));
 sky130_fd_sc_hd__o2111ai_4 _4068_ (.A1(_3243_),
    .A2(_3248_),
    .B1(_3267_),
    .C1(_3268_),
    .D1(_3274_),
    .Y(_3275_));
 sky130_fd_sc_hd__a21oi_1 _4069_ (.A1(_3270_),
    .A2(_3272_),
    .B1(_3273_),
    .Y(_3276_));
 sky130_fd_sc_hd__and3_1 _4070_ (.A(_3269_),
    .B(_3271_),
    .C(_3273_),
    .X(_3277_));
 sky130_fd_sc_hd__o2bb2ai_1 _4071_ (.A1_N(_3268_),
    .A2_N(_3267_),
    .B1(_3276_),
    .B2(_3277_),
    .Y(_3278_));
 sky130_fd_sc_hd__nand4_4 _4072_ (.A(_3205_),
    .B(_3231_),
    .C(_3275_),
    .D(_3278_),
    .Y(_3279_));
 sky130_fd_sc_hd__inv_2 _4073_ (.A(_3279_),
    .Y(_3280_));
 sky130_fd_sc_hd__and3_2 _4074_ (.A(_3210_),
    .B(_3213_),
    .C(_3214_),
    .X(_3281_));
 sky130_fd_sc_hd__a21o_2 _4075_ (.A1(_3222_),
    .A2(_3223_),
    .B1(_3224_),
    .X(_3282_));
 sky130_fd_sc_hd__a31oi_4 _4076_ (.A1(_3216_),
    .A2(_3218_),
    .A3(_3219_),
    .B1(_3282_),
    .Y(_3283_));
 sky130_fd_sc_hd__nand2_1 _4077_ (.A(net285),
    .B(net158),
    .Y(_3284_));
 sky130_fd_sc_hd__nand2_1 _4078_ (.A(net298),
    .B(net152),
    .Y(_3285_));
 sky130_fd_sc_hd__nand2_4 _4079_ (.A(net298),
    .B(net158),
    .Y(_3286_));
 sky130_fd_sc_hd__nand2_4 _4080_ (.A(net285),
    .B(net152),
    .Y(_3287_));
 sky130_fd_sc_hd__o2bb2ai_1 _4081_ (.A1_N(_3284_),
    .A2_N(_3285_),
    .B1(_3286_),
    .B2(_3287_),
    .Y(_3288_));
 sky130_fd_sc_hd__nand3_1 _4082_ (.A(_3288_),
    .B(net163),
    .C(net272),
    .Y(_3289_));
 sky130_fd_sc_hd__nand2_1 _4083_ (.A(net285),
    .B(net165),
    .Y(_3290_));
 sky130_fd_sc_hd__nand2_2 _4084_ (.A(_3286_),
    .B(_3290_),
    .Y(_3291_));
 sky130_fd_sc_hd__nand2_2 _4085_ (.A(net271),
    .B(net174),
    .Y(_3292_));
 sky130_fd_sc_hd__o21ai_1 _4086_ (.A1(_3286_),
    .A2(_3290_),
    .B1(_3292_),
    .Y(_3293_));
 sky130_fd_sc_hd__nand2_1 _4087_ (.A(_3291_),
    .B(_3293_),
    .Y(_3294_));
 sky130_fd_sc_hd__inv_2 _4088_ (.A(net166),
    .Y(_3295_));
 sky130_fd_sc_hd__nand2_2 _4089_ (.A(_3284_),
    .B(_3285_),
    .Y(_3296_));
 sky130_fd_sc_hd__o221ai_4 _4090_ (.A1(_2927_),
    .A2(_3295_),
    .B1(_3287_),
    .B2(_3286_),
    .C1(_3296_),
    .Y(_3297_));
 sky130_fd_sc_hd__nand3_2 _4091_ (.A(_3289_),
    .B(_3294_),
    .C(_3297_),
    .Y(_3298_));
 sky130_fd_sc_hd__and4_1 _4092_ (.A(net298),
    .B(net285),
    .C(net163),
    .D(net156),
    .X(_3299_));
 sky130_fd_sc_hd__a21oi_2 _4093_ (.A1(_3286_),
    .A2(_3290_),
    .B1(_3292_),
    .Y(_3300_));
 sky130_fd_sc_hd__o2111ai_4 _4094_ (.A1(_3287_),
    .A2(_3286_),
    .B1(net271),
    .C1(net165),
    .D1(_3296_),
    .Y(_3301_));
 sky130_fd_sc_hd__o21ai_1 _4095_ (.A1(_2927_),
    .A2(_3295_),
    .B1(_3288_),
    .Y(_3302_));
 sky130_fd_sc_hd__o211ai_4 _4096_ (.A1(_3299_),
    .A2(_3300_),
    .B1(_3301_),
    .C1(_3302_),
    .Y(_3303_));
 sky130_fd_sc_hd__nand4_2 _4097_ (.A(_3298_),
    .B(_3303_),
    .C(net257),
    .D(net170),
    .Y(_3304_));
 sky130_fd_sc_hd__a22o_1 _4098_ (.A1(net256),
    .A2(net170),
    .B1(_3298_),
    .B2(_3303_),
    .X(_3305_));
 sky130_fd_sc_hd__o211ai_4 _4099_ (.A1(_3281_),
    .A2(_3283_),
    .B1(_3304_),
    .C1(_3305_),
    .Y(_3306_));
 sky130_fd_sc_hd__a21oi_1 _4100_ (.A1(_3225_),
    .A2(_3220_),
    .B1(_3281_),
    .Y(_3307_));
 sky130_fd_sc_hd__o211ai_2 _4101_ (.A1(_3176_),
    .A2(_3178_),
    .B1(_3298_),
    .C1(_3303_),
    .Y(_3308_));
 sky130_fd_sc_hd__a21o_1 _4102_ (.A1(_3298_),
    .A2(_3303_),
    .B1(_1147_),
    .X(_3309_));
 sky130_fd_sc_hd__nand3_2 _4103_ (.A(_3307_),
    .B(_3308_),
    .C(_3309_),
    .Y(_3310_));
 sky130_fd_sc_hd__nand4_4 _4104_ (.A(net298),
    .B(net285),
    .C(net165),
    .D(net158),
    .Y(_3311_));
 sky130_fd_sc_hd__a21oi_1 _4105_ (.A1(_3311_),
    .A2(_3291_),
    .B1(_3292_),
    .Y(_3312_));
 sky130_fd_sc_hd__buf_4 _4106_ (.A(_3177_),
    .X(_3313_));
 sky130_fd_sc_hd__o211a_1 _4107_ (.A1(_2927_),
    .A2(_3313_),
    .B1(_3311_),
    .C1(_3291_),
    .X(_3314_));
 sky130_fd_sc_hd__nand4_2 _4108_ (.A(net296),
    .B(net311),
    .C(net169),
    .D(net162),
    .Y(_3315_));
 sky130_fd_sc_hd__nand2_1 _4109_ (.A(net284),
    .B(net174),
    .Y(_3316_));
 sky130_fd_sc_hd__a22oi_4 _4110_ (.A1(net297),
    .A2(net169),
    .B1(net162),
    .B2(net310),
    .Y(_3317_));
 sky130_fd_sc_hd__a21o_2 _4111_ (.A1(_3315_),
    .A2(_3316_),
    .B1(_3317_),
    .X(_3318_));
 sky130_fd_sc_hd__o21bai_4 _4112_ (.A1(_3312_),
    .A2(_3314_),
    .B1_N(_3318_),
    .Y(_3319_));
 sky130_fd_sc_hd__a21oi_1 _4113_ (.A1(_3306_),
    .A2(_3310_),
    .B1(_3319_),
    .Y(_3320_));
 sky130_fd_sc_hd__and3_1 _4114_ (.A(_3319_),
    .B(_3306_),
    .C(_3310_),
    .X(_3321_));
 sky130_fd_sc_hd__a21oi_1 _4115_ (.A1(_3215_),
    .A2(_3221_),
    .B1(_3282_),
    .Y(_3322_));
 sky130_fd_sc_hd__and3_1 _4116_ (.A(_3221_),
    .B(_3282_),
    .C(_3215_),
    .X(_3323_));
 sky130_fd_sc_hd__o21ai_2 _4117_ (.A1(_3322_),
    .A2(_3323_),
    .B1(_3205_),
    .Y(_3324_));
 sky130_fd_sc_hd__a21oi_1 _4118_ (.A1(_3270_),
    .A2(_3272_),
    .B1(_3242_),
    .Y(_3325_));
 sky130_fd_sc_hd__and3_1 _4119_ (.A(_3270_),
    .B(_3272_),
    .C(_3242_),
    .X(_3326_));
 sky130_fd_sc_hd__o2bb2ai_1 _4120_ (.A1_N(_3268_),
    .A2_N(_3267_),
    .B1(_3325_),
    .B2(_3326_),
    .Y(_3327_));
 sky130_fd_sc_hd__a21o_1 _4121_ (.A1(_3270_),
    .A2(_3272_),
    .B1(_3242_),
    .X(_3328_));
 sky130_fd_sc_hd__o22a_2 _4122_ (.A1(_2973_),
    .A2(_3050_),
    .B1(_3207_),
    .B2(_3208_),
    .X(_3329_));
 sky130_fd_sc_hd__o211ai_4 _4123_ (.A1(_3241_),
    .A2(_3329_),
    .B1(_3270_),
    .C1(_3272_),
    .Y(_3330_));
 sky130_fd_sc_hd__nand4_2 _4124_ (.A(_3268_),
    .B(_3267_),
    .C(_3328_),
    .D(_3330_),
    .Y(_3331_));
 sky130_fd_sc_hd__nand4_4 _4125_ (.A(_3230_),
    .B(_3324_),
    .C(_3327_),
    .D(_3331_),
    .Y(_3332_));
 sky130_fd_sc_hd__o211a_1 _4126_ (.A1(_3320_),
    .A2(_3321_),
    .B1(_3332_),
    .C1(_3279_),
    .X(_3333_));
 sky130_fd_sc_hd__and4_1 _4127_ (.A(net298),
    .B(net285),
    .C(net158),
    .D(net152),
    .X(_3334_));
 sky130_fd_sc_hd__nand2_1 _4128_ (.A(net271),
    .B(net165),
    .Y(_3335_));
 sky130_fd_sc_hd__a21oi_2 _4129_ (.A1(_3284_),
    .A2(_3285_),
    .B1(_3335_),
    .Y(_3336_));
 sky130_fd_sc_hd__nand3_2 _4130_ (.A(net256),
    .B(net163),
    .C(net156),
    .Y(_3337_));
 sky130_fd_sc_hd__nand2_1 _4131_ (.A(net256),
    .B(net163),
    .Y(_3338_));
 sky130_fd_sc_hd__nand2_1 _4132_ (.A(net271),
    .B(net156),
    .Y(_3339_));
 sky130_fd_sc_hd__nand2_1 _4133_ (.A(_3338_),
    .B(_3339_),
    .Y(_3340_));
 sky130_fd_sc_hd__o211ai_4 _4134_ (.A1(_2927_),
    .A2(_3337_),
    .B1(_3085_),
    .C1(_3340_),
    .Y(_3341_));
 sky130_fd_sc_hd__clkbuf_8 _4135_ (.A(_1412_),
    .X(_3342_));
 sky130_fd_sc_hd__nand3_1 _4136_ (.A(_3339_),
    .B(net163),
    .C(net256),
    .Y(_3343_));
 sky130_fd_sc_hd__nand3_1 _4137_ (.A(_3338_),
    .B(net156),
    .C(net271),
    .Y(_3344_));
 sky130_fd_sc_hd__o211ai_4 _4138_ (.A1(_3342_),
    .A2(_3313_),
    .B1(_3343_),
    .C1(_3344_),
    .Y(_3345_));
 sky130_fd_sc_hd__o211ai_4 _4139_ (.A1(_3334_),
    .A2(_3336_),
    .B1(_3341_),
    .C1(_3345_),
    .Y(_3346_));
 sky130_fd_sc_hd__o21ai_2 _4140_ (.A1(_3241_),
    .A2(_3329_),
    .B1(_3271_),
    .Y(_3347_));
 sky130_fd_sc_hd__a31o_1 _4141_ (.A1(net271),
    .A2(_3296_),
    .A3(net165),
    .B1(_3334_),
    .X(_3348_));
 sky130_fd_sc_hd__a21o_1 _4142_ (.A1(_3341_),
    .A2(_3345_),
    .B1(_3348_),
    .X(_3349_));
 sky130_fd_sc_hd__nand4_2 _4143_ (.A(_3346_),
    .B(_3270_),
    .C(_3347_),
    .D(_3349_),
    .Y(_3350_));
 sky130_fd_sc_hd__o211a_2 _4144_ (.A1(_3334_),
    .A2(_3336_),
    .B1(_3341_),
    .C1(_3345_),
    .X(_3351_));
 sky130_fd_sc_hd__a21oi_2 _4145_ (.A1(_3341_),
    .A2(_3345_),
    .B1(_3348_),
    .Y(_3352_));
 sky130_fd_sc_hd__o211ai_4 _4146_ (.A1(_3351_),
    .A2(_3352_),
    .B1(_3243_),
    .C1(_3272_),
    .Y(_3353_));
 sky130_fd_sc_hd__nand2_1 _4147_ (.A(_3350_),
    .B(_3353_),
    .Y(_3354_));
 sky130_fd_sc_hd__a32o_1 _4148_ (.A1(_3294_),
    .A2(_3297_),
    .A3(_3289_),
    .B1(_3303_),
    .B2(_1156_),
    .X(_3355_));
 sky130_fd_sc_hd__clkbuf_2 _4149_ (.A(_3355_),
    .X(_3356_));
 sky130_fd_sc_hd__and2_1 _4150_ (.A(_3354_),
    .B(_3356_),
    .X(_3357_));
 sky130_fd_sc_hd__nor2_1 _4151_ (.A(_3354_),
    .B(_3356_),
    .Y(_3358_));
 sky130_fd_sc_hd__o2bb2a_1 _4152_ (.A1_N(_3258_),
    .A2_N(_3264_),
    .B1(_3265_),
    .B2(_3266_),
    .X(_3359_));
 sky130_fd_sc_hd__a31o_1 _4153_ (.A1(_3268_),
    .A2(_3328_),
    .A3(_3330_),
    .B1(_3359_),
    .X(_3360_));
 sky130_fd_sc_hd__o211ai_4 _4154_ (.A1(_3126_),
    .A2(_3127_),
    .B1(_3128_),
    .C1(_3129_),
    .Y(_3361_));
 sky130_fd_sc_hd__nand3_4 _4155_ (.A(_3135_),
    .B(_3132_),
    .C(_3133_),
    .Y(_3362_));
 sky130_fd_sc_hd__o221a_1 _4156_ (.A1(_1793_),
    .A2(_2931_),
    .B1(_2974_),
    .B2(_3093_),
    .C1(_3136_),
    .X(_3363_));
 sky130_fd_sc_hd__o211a_1 _4157_ (.A1(_3095_),
    .A2(_3138_),
    .B1(net322),
    .C1(net135),
    .X(_3364_));
 sky130_fd_sc_hd__o2bb2ai_2 _4158_ (.A1_N(_3361_),
    .A2_N(_3362_),
    .B1(_3363_),
    .B2(_3364_),
    .Y(_3365_));
 sky130_fd_sc_hd__nand4_2 _4159_ (.A(_3361_),
    .B(_3362_),
    .C(_3137_),
    .D(_3139_),
    .Y(_3366_));
 sky130_fd_sc_hd__and4_1 _4160_ (.A(net108),
    .B(net383),
    .C(_3228_),
    .D(_1869_),
    .X(_3367_));
 sky130_fd_sc_hd__a31oi_4 _4161_ (.A1(_3251_),
    .A2(_3254_),
    .A3(_3257_),
    .B1(_3367_),
    .Y(_3368_));
 sky130_fd_sc_hd__nand3_4 _4162_ (.A(_3365_),
    .B(_3366_),
    .C(_3368_),
    .Y(_3369_));
 sky130_fd_sc_hd__a31oi_4 _4163_ (.A1(_3361_),
    .A2(_3362_),
    .A3(_3140_),
    .B1(_3368_),
    .Y(_3370_));
 sky130_fd_sc_hd__a21o_2 _4164_ (.A1(_3361_),
    .A2(_3362_),
    .B1(_3140_),
    .X(_3371_));
 sky130_fd_sc_hd__nand2_4 _4165_ (.A(_3370_),
    .B(_3371_),
    .Y(_3372_));
 sky130_fd_sc_hd__nand4_1 _4166_ (.A(net297),
    .B(net310),
    .C(net146),
    .D(net140),
    .Y(_3373_));
 sky130_fd_sc_hd__a22oi_1 _4167_ (.A1(net283),
    .A2(net151),
    .B1(_3103_),
    .B2(_3373_),
    .Y(_3374_));
 sky130_fd_sc_hd__o21ai_1 _4168_ (.A1(_3092_),
    .A2(_3252_),
    .B1(_3256_),
    .Y(_3375_));
 sky130_fd_sc_hd__o2111ai_1 _4169_ (.A1(_1231_),
    .A2(_3237_),
    .B1(net284),
    .C1(net151),
    .D1(_3103_),
    .Y(_3376_));
 sky130_fd_sc_hd__nand3b_1 _4170_ (.A_N(_3374_),
    .B(_3375_),
    .C(_3376_),
    .Y(_3377_));
 sky130_fd_sc_hd__buf_2 _4171_ (.A(_3377_),
    .X(_3378_));
 sky130_fd_sc_hd__o22a_1 _4172_ (.A1(_2981_),
    .A2(_3182_),
    .B1(_3092_),
    .B2(_3252_),
    .X(_3379_));
 sky130_fd_sc_hd__a21o_1 _4173_ (.A1(_3103_),
    .A2(_3373_),
    .B1(_3287_),
    .X(_3380_));
 sky130_fd_sc_hd__inv_6 _4174_ (.A(net284),
    .Y(_3381_));
 sky130_fd_sc_hd__o221ai_2 _4175_ (.A1(_3381_),
    .A2(_1445_),
    .B1(_1231_),
    .B2(_3237_),
    .C1(_3103_),
    .Y(_3382_));
 sky130_fd_sc_hd__nand3_1 _4176_ (.A(_3379_),
    .B(_3380_),
    .C(_3382_),
    .Y(_3383_));
 sky130_fd_sc_hd__clkbuf_2 _4177_ (.A(_3383_),
    .X(_3384_));
 sky130_fd_sc_hd__o32a_2 _4178_ (.A1(_1793_),
    .A2(_2931_),
    .A3(_3207_),
    .B1(_3245_),
    .B2(_3237_),
    .X(_3385_));
 sky130_fd_sc_hd__a21oi_1 _4179_ (.A1(_3378_),
    .A2(_3384_),
    .B1(_3385_),
    .Y(_3386_));
 sky130_fd_sc_hd__and3_1 _4180_ (.A(_3378_),
    .B(_3384_),
    .C(_3385_),
    .X(_3387_));
 sky130_fd_sc_hd__o2bb2ai_2 _4181_ (.A1_N(_3369_),
    .A2_N(_3372_),
    .B1(_3386_),
    .B2(_3387_),
    .Y(_3388_));
 sky130_fd_sc_hd__a21boi_2 _4182_ (.A1(_3378_),
    .A2(_3384_),
    .B1_N(_3385_),
    .Y(_3389_));
 sky130_fd_sc_hd__and3b_1 _4183_ (.A_N(_3385_),
    .B(_3384_),
    .C(_3378_),
    .X(_3390_));
 sky130_fd_sc_hd__o211ai_4 _4184_ (.A1(_3389_),
    .A2(_3390_),
    .B1(_3369_),
    .C1(_3372_),
    .Y(_3391_));
 sky130_fd_sc_hd__o2111ai_2 _4185_ (.A1(_3357_),
    .A2(_3358_),
    .B1(_3360_),
    .C1(_3388_),
    .D1(_3391_),
    .Y(_3392_));
 sky130_fd_sc_hd__a31oi_2 _4186_ (.A1(_3268_),
    .A2(_3328_),
    .A3(_3330_),
    .B1(_3359_),
    .Y(_3393_));
 sky130_fd_sc_hd__o211ai_2 _4187_ (.A1(_3386_),
    .A2(_3387_),
    .B1(_3369_),
    .C1(_3372_),
    .Y(_3394_));
 sky130_fd_sc_hd__nand2_1 _4188_ (.A(_3354_),
    .B(_3356_),
    .Y(_3395_));
 sky130_fd_sc_hd__nand3b_1 _4189_ (.A_N(_3355_),
    .B(_3353_),
    .C(_3350_),
    .Y(_3396_));
 sky130_fd_sc_hd__nand4_1 _4190_ (.A(_3393_),
    .B(_3394_),
    .C(_3395_),
    .D(_3396_),
    .Y(_3397_));
 sky130_fd_sc_hd__a21o_1 _4191_ (.A1(_3377_),
    .A2(_3383_),
    .B1(_3385_),
    .X(_3398_));
 sky130_fd_sc_hd__o2111ai_1 _4192_ (.A1(_3237_),
    .A2(_3245_),
    .B1(_3235_),
    .C1(_3378_),
    .D1(_3384_),
    .Y(_3399_));
 sky130_fd_sc_hd__nand2_1 _4193_ (.A(_3398_),
    .B(_3399_),
    .Y(_3400_));
 sky130_fd_sc_hd__a21oi_2 _4194_ (.A1(_3369_),
    .A2(_3372_),
    .B1(_3400_),
    .Y(_3401_));
 sky130_fd_sc_hd__nand3_2 _4195_ (.A(_3388_),
    .B(_3391_),
    .C(_3360_),
    .Y(_3402_));
 sky130_fd_sc_hd__nand2_1 _4196_ (.A(_3393_),
    .B(_3394_),
    .Y(_3403_));
 sky130_fd_sc_hd__nand2_1 _4197_ (.A(_3395_),
    .B(_3396_),
    .Y(_3404_));
 sky130_fd_sc_hd__o21ai_1 _4198_ (.A1(_3401_),
    .A2(_3403_),
    .B1(_3404_),
    .Y(_3405_));
 sky130_fd_sc_hd__o211ai_2 _4199_ (.A1(_3397_),
    .A2(_3401_),
    .B1(_3402_),
    .C1(_3405_),
    .Y(_3406_));
 sky130_fd_sc_hd__o211ai_1 _4200_ (.A1(_3280_),
    .A2(_3333_),
    .B1(_3392_),
    .C1(_3406_),
    .Y(_3407_));
 sky130_fd_sc_hd__inv_2 _4201_ (.A(_3402_),
    .Y(_3408_));
 sky130_fd_sc_hd__a21o_1 _4202_ (.A1(_3311_),
    .A2(_3291_),
    .B1(_3292_),
    .X(_3409_));
 sky130_fd_sc_hd__o211ai_4 _4203_ (.A1(_2928_),
    .A2(_3178_),
    .B1(_3311_),
    .C1(_3291_),
    .Y(_3410_));
 sky130_fd_sc_hd__a21oi_2 _4204_ (.A1(_3409_),
    .A2(_3410_),
    .B1(_3318_),
    .Y(_3411_));
 sky130_fd_sc_hd__a21o_1 _4205_ (.A1(_3306_),
    .A2(_3310_),
    .B1(_3411_),
    .X(_3412_));
 sky130_fd_sc_hd__nand3_2 _4206_ (.A(_3306_),
    .B(_3310_),
    .C(_3411_),
    .Y(_3413_));
 sky130_fd_sc_hd__a31oi_2 _4207_ (.A1(_3332_),
    .A2(_3412_),
    .A3(_3413_),
    .B1(_3280_),
    .Y(_3414_));
 sky130_fd_sc_hd__o2bb2ai_1 _4208_ (.A1_N(_3369_),
    .A2_N(_3372_),
    .B1(_3389_),
    .B2(_3390_),
    .Y(_3415_));
 sky130_fd_sc_hd__nand3_1 _4209_ (.A(_3393_),
    .B(_3415_),
    .C(_3394_),
    .Y(_3416_));
 sky130_fd_sc_hd__a21oi_1 _4210_ (.A1(_3350_),
    .A2(_3353_),
    .B1(_3356_),
    .Y(_3417_));
 sky130_fd_sc_hd__and3_1 _4211_ (.A(_3350_),
    .B(_3353_),
    .C(_3356_),
    .X(_3418_));
 sky130_fd_sc_hd__o2bb2ai_1 _4212_ (.A1_N(_3402_),
    .A2_N(_3416_),
    .B1(_3417_),
    .B2(_3418_),
    .Y(_3419_));
 sky130_fd_sc_hd__o211ai_1 _4213_ (.A1(_3405_),
    .A2(_3408_),
    .B1(_3414_),
    .C1(_3419_),
    .Y(_3420_));
 sky130_fd_sc_hd__inv_2 _4214_ (.A(_3306_),
    .Y(_3421_));
 sky130_fd_sc_hd__a21o_1 _4215_ (.A1(_3411_),
    .A2(_3310_),
    .B1(_3421_),
    .X(_3422_));
 sky130_fd_sc_hd__a21o_1 _4216_ (.A1(_3407_),
    .A2(_3420_),
    .B1(_3422_),
    .X(_3423_));
 sky130_fd_sc_hd__o22a_1 _4217_ (.A1(_3357_),
    .A2(_3358_),
    .B1(_3401_),
    .B2(_3403_),
    .X(_3424_));
 sky130_fd_sc_hd__nand2_1 _4218_ (.A(_3424_),
    .B(_3402_),
    .Y(_3425_));
 sky130_fd_sc_hd__a21oi_1 _4219_ (.A1(_3411_),
    .A2(_3310_),
    .B1(_3421_),
    .Y(_3426_));
 sky130_fd_sc_hd__a31oi_2 _4220_ (.A1(_3425_),
    .A2(_3419_),
    .A3(_3414_),
    .B1(_3426_),
    .Y(_3427_));
 sky130_fd_sc_hd__nand2_1 _4221_ (.A(_3427_),
    .B(_3407_),
    .Y(_3428_));
 sky130_fd_sc_hd__nand3_4 _4222_ (.A(_3409_),
    .B(_3410_),
    .C(_3318_),
    .Y(_3429_));
 sky130_fd_sc_hd__nand2_1 _4223_ (.A(net374),
    .B(net134),
    .Y(_3430_));
 sky130_fd_sc_hd__a22oi_4 _4224_ (.A1(net120),
    .A2(net394),
    .B1(net384),
    .B2(net126),
    .Y(_3431_));
 sky130_fd_sc_hd__nand4_2 _4225_ (.A(net120),
    .B(net395),
    .C(net384),
    .D(net126),
    .Y(_3432_));
 sky130_fd_sc_hd__o21a_1 _4226_ (.A1(_3430_),
    .A2(_3431_),
    .B1(_3432_),
    .X(_3433_));
 sky130_fd_sc_hd__nand2_2 _4227_ (.A(net350),
    .B(net142),
    .Y(_3434_));
 sky130_fd_sc_hd__nand2_1 _4228_ (.A(net336),
    .B(net146),
    .Y(_3435_));
 sky130_fd_sc_hd__nand2_2 _4229_ (.A(_3434_),
    .B(_3435_),
    .Y(_3436_));
 sky130_fd_sc_hd__a21o_1 _4230_ (.A1(_3436_),
    .A2(_3223_),
    .B1(_3222_),
    .X(_3437_));
 sky130_fd_sc_hd__o211ai_2 _4231_ (.A1(_2886_),
    .A2(_1445_),
    .B1(_3436_),
    .C1(_3223_),
    .Y(_3438_));
 sky130_fd_sc_hd__nand3_4 _4232_ (.A(_3433_),
    .B(_3437_),
    .C(_3438_),
    .Y(_3439_));
 sky130_fd_sc_hd__a22oi_4 _4233_ (.A1(net349),
    .A2(net147),
    .B1(net139),
    .B2(net361),
    .Y(_3440_));
 sky130_fd_sc_hd__buf_6 _4234_ (.A(_2120_),
    .X(_3441_));
 sky130_fd_sc_hd__nand2_2 _4235_ (.A(net359),
    .B(net148),
    .Y(_3442_));
 sky130_fd_sc_hd__o22a_2 _4236_ (.A1(_3441_),
    .A2(_3050_),
    .B1(_3434_),
    .B2(_3442_),
    .X(_3443_));
 sky130_fd_sc_hd__o2bb2ai_2 _4237_ (.A1_N(_3436_),
    .A2_N(_3223_),
    .B1(_1782_),
    .B2(_1445_),
    .Y(_3444_));
 sky130_fd_sc_hd__nand4_2 _4238_ (.A(_3436_),
    .B(_3223_),
    .C(net323),
    .D(net153),
    .Y(_3445_));
 sky130_fd_sc_hd__o21ai_2 _4239_ (.A1(_3430_),
    .A2(_3431_),
    .B1(_3432_),
    .Y(_3446_));
 sky130_fd_sc_hd__nand3_4 _4240_ (.A(_3444_),
    .B(_3445_),
    .C(_3446_),
    .Y(_3447_));
 sky130_fd_sc_hd__o21ai_1 _4241_ (.A1(_3440_),
    .A2(_3443_),
    .B1(_3447_),
    .Y(_3448_));
 sky130_fd_sc_hd__nand4_4 _4242_ (.A(_3319_),
    .B(_3429_),
    .C(_3439_),
    .D(_3448_),
    .Y(_3449_));
 sky130_fd_sc_hd__nand2_2 _4243_ (.A(net325),
    .B(net161),
    .Y(_3450_));
 sky130_fd_sc_hd__nand2_1 _4244_ (.A(net314),
    .B(net166),
    .Y(_3451_));
 sky130_fd_sc_hd__nand2_2 _4245_ (.A(_3450_),
    .B(_3451_),
    .Y(_3452_));
 sky130_fd_sc_hd__nand2_1 _4246_ (.A(net304),
    .B(net173),
    .Y(_3453_));
 sky130_fd_sc_hd__o21ai_1 _4247_ (.A1(_3450_),
    .A2(_3451_),
    .B1(_3453_),
    .Y(_3454_));
 sky130_fd_sc_hd__nand2_2 _4248_ (.A(_3452_),
    .B(_3454_),
    .Y(_3455_));
 sky130_fd_sc_hd__and4_1 _4249_ (.A(net297),
    .B(net310),
    .C(net169),
    .D(net162),
    .X(_3456_));
 sky130_fd_sc_hd__o21ai_1 _4250_ (.A1(_3456_),
    .A2(_3317_),
    .B1(_3316_),
    .Y(_3457_));
 sky130_fd_sc_hd__nand4b_1 _4251_ (.A_N(_3317_),
    .B(net174),
    .C(net284),
    .D(_3315_),
    .Y(_3458_));
 sky130_fd_sc_hd__nand3b_2 _4252_ (.A_N(_3455_),
    .B(_3457_),
    .C(_3458_),
    .Y(_3459_));
 sky130_fd_sc_hd__a21oi_1 _4253_ (.A1(_3444_),
    .A2(_3445_),
    .B1(_3446_),
    .Y(_3460_));
 sky130_fd_sc_hd__nand4_1 _4254_ (.A(net361),
    .B(net349),
    .C(net146),
    .D(net142),
    .Y(_3461_));
 sky130_fd_sc_hd__o31a_1 _4255_ (.A1(_3441_),
    .A2(_3050_),
    .A3(_3440_),
    .B1(_3461_),
    .X(_3462_));
 sky130_fd_sc_hd__nand2_1 _4256_ (.A(_3319_),
    .B(_3429_),
    .Y(_3463_));
 sky130_fd_sc_hd__o211ai_2 _4257_ (.A1(_3460_),
    .A2(_3462_),
    .B1(_3447_),
    .C1(_3463_),
    .Y(_3464_));
 sky130_fd_sc_hd__nand3b_2 _4258_ (.A_N(_3459_),
    .B(_3464_),
    .C(_3449_),
    .Y(_3465_));
 sky130_fd_sc_hd__and2_1 _4259_ (.A(_3449_),
    .B(_3465_),
    .X(_3466_));
 sky130_fd_sc_hd__inv_2 _4260_ (.A(_3466_),
    .Y(_3467_));
 sky130_fd_sc_hd__a21oi_1 _4261_ (.A1(_3306_),
    .A2(_3310_),
    .B1(_3411_),
    .Y(_3468_));
 sky130_fd_sc_hd__inv_2 _4262_ (.A(_3413_),
    .Y(_3469_));
 sky130_fd_sc_hd__o211ai_1 _4263_ (.A1(_3468_),
    .A2(_3469_),
    .B1(_3332_),
    .C1(_3279_),
    .Y(_3470_));
 sky130_fd_sc_hd__o2bb2ai_1 _4264_ (.A1_N(_3332_),
    .A2_N(_3279_),
    .B1(_3320_),
    .B2(_3321_),
    .Y(_3471_));
 sky130_fd_sc_hd__a21oi_2 _4265_ (.A1(_3201_),
    .A2(_3202_),
    .B1(_3204_),
    .Y(_3472_));
 sky130_fd_sc_hd__and3_1 _4266_ (.A(_3204_),
    .B(_3201_),
    .C(_3202_),
    .X(_3473_));
 sky130_fd_sc_hd__and4_1 _4267_ (.A(net361),
    .B(net350),
    .C(net147),
    .D(net142),
    .X(_3474_));
 sky130_fd_sc_hd__and2_1 _4268_ (.A(net336),
    .B(net153),
    .X(_3475_));
 sky130_fd_sc_hd__nand2_1 _4269_ (.A(net347),
    .B(net146),
    .Y(_3476_));
 sky130_fd_sc_hd__nand2_1 _4270_ (.A(net361),
    .B(net141),
    .Y(_3477_));
 sky130_fd_sc_hd__nand2_4 _4271_ (.A(_3476_),
    .B(_3477_),
    .Y(_3478_));
 sky130_fd_sc_hd__o2111ai_4 _4272_ (.A1(_3474_),
    .A2(_3475_),
    .B1(_3478_),
    .C1(_3439_),
    .D1(_3447_),
    .Y(_3479_));
 sky130_fd_sc_hd__o2bb2ai_1 _4273_ (.A1_N(_3439_),
    .A2_N(_3447_),
    .B1(_3440_),
    .B2(_3443_),
    .Y(_3480_));
 sky130_fd_sc_hd__o211ai_4 _4274_ (.A1(_3472_),
    .A2(_3473_),
    .B1(_3479_),
    .C1(_3480_),
    .Y(_3481_));
 sky130_fd_sc_hd__a21o_1 _4275_ (.A1(_3215_),
    .A2(_3221_),
    .B1(_3282_),
    .X(_3482_));
 sky130_fd_sc_hd__nand3_1 _4276_ (.A(_3221_),
    .B(_3282_),
    .C(_3215_),
    .Y(_3483_));
 sky130_fd_sc_hd__nand4_1 _4277_ (.A(_3205_),
    .B(_3230_),
    .C(_3482_),
    .D(_3483_),
    .Y(_3484_));
 sky130_fd_sc_hd__o2bb2ai_1 _4278_ (.A1_N(_3205_),
    .A2_N(_3230_),
    .B1(_3322_),
    .B2(_3323_),
    .Y(_3485_));
 sky130_fd_sc_hd__nand3_2 _4279_ (.A(_3481_),
    .B(_3484_),
    .C(_3485_),
    .Y(_3486_));
 sky130_fd_sc_hd__o21ai_2 _4280_ (.A1(_3381_),
    .A2(_3313_),
    .B1(_3315_),
    .Y(_3487_));
 sky130_fd_sc_hd__o21bai_2 _4281_ (.A1(_3456_),
    .A2(_3317_),
    .B1_N(_3316_),
    .Y(_3488_));
 sky130_fd_sc_hd__o21a_1 _4282_ (.A1(_3317_),
    .A2(_3487_),
    .B1(_3488_),
    .X(_3489_));
 sky130_fd_sc_hd__o2bb2ai_2 _4283_ (.A1_N(_3449_),
    .A2_N(_3464_),
    .B1(_3489_),
    .B2(_3455_),
    .Y(_3490_));
 sky130_fd_sc_hd__a21oi_1 _4284_ (.A1(_3484_),
    .A2(_3485_),
    .B1(_3481_),
    .Y(_3491_));
 sky130_fd_sc_hd__a31oi_2 _4285_ (.A1(_3465_),
    .A2(_3486_),
    .A3(_3490_),
    .B1(_3491_),
    .Y(_3492_));
 sky130_fd_sc_hd__nand3_2 _4286_ (.A(_3470_),
    .B(_3471_),
    .C(_3492_),
    .Y(_3493_));
 sky130_fd_sc_hd__nand4_1 _4287_ (.A(_3332_),
    .B(_3279_),
    .C(_3412_),
    .D(_3413_),
    .Y(_3494_));
 sky130_fd_sc_hd__o2bb2ai_1 _4288_ (.A1_N(_3332_),
    .A2_N(_3279_),
    .B1(_3468_),
    .B2(_3469_),
    .Y(_3495_));
 sky130_fd_sc_hd__a31o_1 _4289_ (.A1(_3216_),
    .A2(_3218_),
    .A3(_3219_),
    .B1(_3282_),
    .X(_3496_));
 sky130_fd_sc_hd__a21o_1 _4290_ (.A1(_3215_),
    .A2(_3221_),
    .B1(_3225_),
    .X(_3497_));
 sky130_fd_sc_hd__o2111ai_2 _4291_ (.A1(_3496_),
    .A2(_3281_),
    .B1(_3230_),
    .C1(_3205_),
    .D1(_3497_),
    .Y(_3498_));
 sky130_fd_sc_hd__o2bb2ai_1 _4292_ (.A1_N(_3205_),
    .A2_N(_3230_),
    .B1(_3226_),
    .B2(_3227_),
    .Y(_3499_));
 sky130_fd_sc_hd__nand3b_2 _4293_ (.A_N(_3481_),
    .B(_3498_),
    .C(_3499_),
    .Y(_3500_));
 sky130_fd_sc_hd__nand2_1 _4294_ (.A(_3465_),
    .B(_3490_),
    .Y(_3501_));
 sky130_fd_sc_hd__a21boi_2 _4295_ (.A1(_3500_),
    .A2(_3501_),
    .B1_N(_3486_),
    .Y(_3502_));
 sky130_fd_sc_hd__nand3_2 _4296_ (.A(_3494_),
    .B(_3495_),
    .C(_3502_),
    .Y(_3503_));
 sky130_fd_sc_hd__a21bo_1 _4297_ (.A1(_3467_),
    .A2(_3493_),
    .B1_N(_3503_),
    .X(_3504_));
 sky130_fd_sc_hd__a21o_1 _4298_ (.A1(_3423_),
    .A2(_3428_),
    .B1(_3504_),
    .X(_3505_));
 sky130_fd_sc_hd__nand3_2 _4299_ (.A(_3423_),
    .B(_3428_),
    .C(_3504_),
    .Y(_3506_));
 sky130_fd_sc_hd__inv_2 _4300_ (.A(_3353_),
    .Y(_3507_));
 sky130_fd_sc_hd__and2_1 _4301_ (.A(_3350_),
    .B(_3356_),
    .X(_3508_));
 sky130_fd_sc_hd__and4_1 _4302_ (.A(net257),
    .B(net174),
    .C(net165),
    .D(net158),
    .X(_3509_));
 sky130_fd_sc_hd__and4_1 _4303_ (.A(net271),
    .B(net257),
    .C(net164),
    .D(net156),
    .X(_3510_));
 sky130_fd_sc_hd__a21oi_1 _4304_ (.A1(_3084_),
    .A2(_3337_),
    .B1(_1147_),
    .Y(_3511_));
 sky130_fd_sc_hd__and3_1 _4305_ (.A(net256),
    .B(net163),
    .C(net157),
    .X(_3512_));
 sky130_fd_sc_hd__o31ai_1 _4306_ (.A1(_3086_),
    .A2(_1174_),
    .A3(_3512_),
    .B1(_3341_),
    .Y(_3513_));
 sky130_fd_sc_hd__nor3_1 _4307_ (.A(_3510_),
    .B(_3511_),
    .C(_3513_),
    .Y(_3514_));
 sky130_fd_sc_hd__a31o_1 _4308_ (.A1(_3379_),
    .A2(_3380_),
    .A3(_3382_),
    .B1(_3385_),
    .X(_3515_));
 sky130_fd_sc_hd__o211ai_4 _4309_ (.A1(_3509_),
    .A2(_3514_),
    .B1(_3515_),
    .C1(_3378_),
    .Y(_3516_));
 sky130_fd_sc_hd__or4b_1 _4310_ (.A(_3342_),
    .B(_3178_),
    .C(_3295_),
    .D_N(net156),
    .X(_3517_));
 sky130_fd_sc_hd__o31a_1 _4311_ (.A1(_3510_),
    .A2(_3511_),
    .A3(_3513_),
    .B1(_3517_),
    .X(_3518_));
 sky130_fd_sc_hd__nand2_1 _4312_ (.A(_3378_),
    .B(_3385_),
    .Y(_3519_));
 sky130_fd_sc_hd__nand3_2 _4313_ (.A(_3518_),
    .B(_3519_),
    .C(_3384_),
    .Y(_3520_));
 sky130_fd_sc_hd__and3_1 _4314_ (.A(_3516_),
    .B(_3520_),
    .C(_3351_),
    .X(_3521_));
 sky130_fd_sc_hd__a21oi_1 _4315_ (.A1(_3516_),
    .A2(_3520_),
    .B1(_3351_),
    .Y(_3522_));
 sky130_fd_sc_hd__o211ai_4 _4316_ (.A1(_3149_),
    .A2(_3154_),
    .B1(_3147_),
    .C1(_3155_),
    .Y(_3523_));
 sky130_fd_sc_hd__nand2_1 _4317_ (.A(_3146_),
    .B(_3523_),
    .Y(_3524_));
 sky130_fd_sc_hd__o21ai_2 _4318_ (.A1(_3121_),
    .A2(_3122_),
    .B1(_3524_),
    .Y(_3525_));
 sky130_fd_sc_hd__a22o_1 _4319_ (.A1(_3370_),
    .A2(_3371_),
    .B1(_3369_),
    .B2(_3400_),
    .X(_3526_));
 sky130_fd_sc_hd__o211ai_2 _4320_ (.A1(_3148_),
    .A2(_3156_),
    .B1(_3123_),
    .C1(_3146_),
    .Y(_3527_));
 sky130_fd_sc_hd__nand3_2 _4321_ (.A(_3525_),
    .B(_3526_),
    .C(_3527_),
    .Y(_3528_));
 sky130_fd_sc_hd__o21ai_1 _4322_ (.A1(_3121_),
    .A2(_3122_),
    .B1(_3146_),
    .Y(_3529_));
 sky130_fd_sc_hd__inv_2 _4323_ (.A(_3523_),
    .Y(_3530_));
 sky130_fd_sc_hd__a22oi_2 _4324_ (.A1(_3370_),
    .A2(_3371_),
    .B1(_3369_),
    .B2(_3400_),
    .Y(_3531_));
 sky130_fd_sc_hd__nand2_1 _4325_ (.A(_3524_),
    .B(_3123_),
    .Y(_3532_));
 sky130_fd_sc_hd__o211ai_4 _4326_ (.A1(_3529_),
    .A2(_3530_),
    .B1(_3531_),
    .C1(_3532_),
    .Y(_3533_));
 sky130_fd_sc_hd__o211ai_2 _4327_ (.A1(_3521_),
    .A2(_3522_),
    .B1(_3528_),
    .C1(_3533_),
    .Y(_3534_));
 sky130_fd_sc_hd__a21oi_1 _4328_ (.A1(_3516_),
    .A2(_3520_),
    .B1(_3346_),
    .Y(_3535_));
 sky130_fd_sc_hd__and3_1 _4329_ (.A(_3346_),
    .B(_3516_),
    .C(_3520_),
    .X(_3536_));
 sky130_fd_sc_hd__o2bb2ai_1 _4330_ (.A1_N(_3528_),
    .A2_N(_3533_),
    .B1(_3535_),
    .B2(_3536_),
    .Y(_3537_));
 sky130_fd_sc_hd__o211ai_4 _4331_ (.A1(_3408_),
    .A2(_3424_),
    .B1(_3534_),
    .C1(_3537_),
    .Y(_0105_));
 sky130_fd_sc_hd__nor2_1 _4332_ (.A(_3521_),
    .B(_3522_),
    .Y(_0106_));
 sky130_fd_sc_hd__a21o_1 _4333_ (.A1(_3528_),
    .A2(_3533_),
    .B1(_0106_),
    .X(_0107_));
 sky130_fd_sc_hd__a32oi_2 _4334_ (.A1(_3360_),
    .A2(_3388_),
    .A3(_3391_),
    .B1(_3416_),
    .B2(_3404_),
    .Y(_0108_));
 sky130_fd_sc_hd__o211ai_1 _4335_ (.A1(_3535_),
    .A2(_3536_),
    .B1(_3528_),
    .C1(_3533_),
    .Y(_0109_));
 sky130_fd_sc_hd__nand3_2 _4336_ (.A(_0107_),
    .B(_0108_),
    .C(_0109_),
    .Y(_0110_));
 sky130_fd_sc_hd__o211a_1 _4337_ (.A1(_3507_),
    .A2(_3508_),
    .B1(_0105_),
    .C1(_0110_),
    .X(_0111_));
 sky130_fd_sc_hd__a21o_1 _4338_ (.A1(_3350_),
    .A2(_3356_),
    .B1(_3507_),
    .X(_0112_));
 sky130_fd_sc_hd__a21o_1 _4339_ (.A1(_0110_),
    .A2(_0105_),
    .B1(_0112_),
    .X(_0113_));
 sky130_fd_sc_hd__o211a_1 _4340_ (.A1(_3280_),
    .A2(_3333_),
    .B1(_3392_),
    .C1(_3406_),
    .X(_0114_));
 sky130_fd_sc_hd__a21oi_1 _4341_ (.A1(_3420_),
    .A2(_3422_),
    .B1(_0114_),
    .Y(_0115_));
 sky130_fd_sc_hd__nand3b_2 _4342_ (.A_N(_0111_),
    .B(_0113_),
    .C(_0115_),
    .Y(_0116_));
 sky130_fd_sc_hd__nand3b_1 _4343_ (.A_N(_0112_),
    .B(_0105_),
    .C(_0110_),
    .Y(_0117_));
 sky130_fd_sc_hd__o2bb2ai_1 _4344_ (.A1_N(_0110_),
    .A2_N(_0105_),
    .B1(_3508_),
    .B2(_3507_),
    .Y(_0118_));
 sky130_fd_sc_hd__o211ai_2 _4345_ (.A1(_0114_),
    .A2(_3427_),
    .B1(_0117_),
    .C1(_0118_),
    .Y(_0119_));
 sky130_fd_sc_hd__nand4_2 _4346_ (.A(_3505_),
    .B(_3506_),
    .C(_0116_),
    .D(_0119_),
    .Y(_0120_));
 sky130_fd_sc_hd__a22o_1 _4347_ (.A1(_3449_),
    .A2(_3465_),
    .B1(_3493_),
    .B2(_3503_),
    .X(_0121_));
 sky130_fd_sc_hd__nand4_1 _4348_ (.A(_3449_),
    .B(_3465_),
    .C(_3493_),
    .D(_3503_),
    .Y(_0122_));
 sky130_fd_sc_hd__and3_1 _4349_ (.A(_3461_),
    .B(_3478_),
    .C(_3475_),
    .X(_0123_));
 sky130_fd_sc_hd__o2bb2ai_1 _4350_ (.A1_N(_3461_),
    .A2_N(_3478_),
    .B1(_2120_),
    .B2(_1445_),
    .Y(_0124_));
 sky130_fd_sc_hd__and4_2 _4351_ (.A(net394),
    .B(net385),
    .C(net135),
    .D(net127),
    .X(_0125_));
 sky130_fd_sc_hd__nand2_1 _4352_ (.A(_0124_),
    .B(_0125_),
    .Y(_0126_));
 sky130_fd_sc_hd__nand4_2 _4353_ (.A(net394),
    .B(net385),
    .C(net135),
    .D(net127),
    .Y(_0127_));
 sky130_fd_sc_hd__o221ai_4 _4354_ (.A1(_2120_),
    .A2(_3049_),
    .B1(_3434_),
    .B2(_3442_),
    .C1(_3478_),
    .Y(_0128_));
 sky130_fd_sc_hd__o21ai_1 _4355_ (.A1(_3434_),
    .A2(_3442_),
    .B1(_3478_),
    .Y(_0129_));
 sky130_fd_sc_hd__nand2_1 _4356_ (.A(_0129_),
    .B(_3475_),
    .Y(_0130_));
 sky130_fd_sc_hd__nand3_4 _4357_ (.A(_0127_),
    .B(_0128_),
    .C(_0130_),
    .Y(_0131_));
 sky130_fd_sc_hd__o21ai_1 _4358_ (.A1(_0123_),
    .A2(_0126_),
    .B1(_0131_),
    .Y(_0132_));
 sky130_fd_sc_hd__nand2_4 _4359_ (.A(net371),
    .B(net359),
    .Y(_0133_));
 sky130_fd_sc_hd__nand2_1 _4360_ (.A(net347),
    .B(net154),
    .Y(_0134_));
 sky130_fd_sc_hd__a22oi_4 _4361_ (.A1(net364),
    .A2(net148),
    .B1(net141),
    .B2(net372),
    .Y(_0135_));
 sky130_fd_sc_hd__o22a_2 _4362_ (.A1(_2555_),
    .A2(_0133_),
    .B1(_0134_),
    .B2(_0135_),
    .X(_0136_));
 sky130_fd_sc_hd__nand2_2 _4363_ (.A(_0132_),
    .B(_0136_),
    .Y(_0137_));
 sky130_fd_sc_hd__a41o_1 _4364_ (.A1(net120),
    .A2(net394),
    .A3(net384),
    .A4(net126),
    .B1(_3430_),
    .X(_0138_));
 sky130_fd_sc_hd__a22o_1 _4365_ (.A1(net120),
    .A2(net394),
    .B1(net384),
    .B2(net126),
    .X(_0139_));
 sky130_fd_sc_hd__a22o_1 _4366_ (.A1(net374),
    .A2(net134),
    .B1(_0139_),
    .B2(_3432_),
    .X(_0140_));
 sky130_fd_sc_hd__o21a_2 _4367_ (.A1(_3431_),
    .A2(_0138_),
    .B1(_0140_),
    .X(_0141_));
 sky130_fd_sc_hd__o2111ai_1 _4368_ (.A1(_3434_),
    .A2(_3442_),
    .B1(net336),
    .C1(net153),
    .D1(_3478_),
    .Y(_0142_));
 sky130_fd_sc_hd__nand3_2 _4369_ (.A(_0124_),
    .B(_0125_),
    .C(_0142_),
    .Y(_0143_));
 sky130_fd_sc_hd__nand3b_4 _4370_ (.A_N(_0136_),
    .B(_0143_),
    .C(_0131_),
    .Y(_0144_));
 sky130_fd_sc_hd__nand3_4 _4371_ (.A(_0137_),
    .B(_0141_),
    .C(_0144_),
    .Y(_0145_));
 sky130_fd_sc_hd__nor2_1 _4372_ (.A(_3472_),
    .B(_3473_),
    .Y(_0146_));
 sky130_fd_sc_hd__a21o_1 _4373_ (.A1(_3439_),
    .A2(_3447_),
    .B1(_3462_),
    .X(_0147_));
 sky130_fd_sc_hd__o211ai_1 _4374_ (.A1(_3440_),
    .A2(_3443_),
    .B1(_3439_),
    .C1(_3447_),
    .Y(_0148_));
 sky130_fd_sc_hd__nand3_2 _4375_ (.A(_0146_),
    .B(_0147_),
    .C(_0148_),
    .Y(_0149_));
 sky130_fd_sc_hd__nand3b_4 _4376_ (.A_N(_0145_),
    .B(_0149_),
    .C(_3481_),
    .Y(_0150_));
 sky130_fd_sc_hd__nand2_1 _4377_ (.A(_0144_),
    .B(_0137_),
    .Y(_0151_));
 sky130_fd_sc_hd__o21ai_1 _4378_ (.A1(_3431_),
    .A2(_0138_),
    .B1(_0140_),
    .Y(_0152_));
 sky130_fd_sc_hd__o2bb2ai_2 _4379_ (.A1_N(_3481_),
    .A2_N(_0149_),
    .B1(_0151_),
    .B2(_0152_),
    .Y(_0153_));
 sky130_fd_sc_hd__o211ai_4 _4380_ (.A1(_3317_),
    .A2(_3487_),
    .B1(_3455_),
    .C1(_3488_),
    .Y(_0154_));
 sky130_fd_sc_hd__nand2_1 _4381_ (.A(_0143_),
    .B(_0136_),
    .Y(_0155_));
 sky130_fd_sc_hd__nand4_4 _4382_ (.A(_3459_),
    .B(_0131_),
    .C(_0154_),
    .D(_0155_),
    .Y(_0156_));
 sky130_fd_sc_hd__a31o_1 _4383_ (.A1(_0127_),
    .A2(_0128_),
    .A3(_0130_),
    .B1(_0136_),
    .X(_0157_));
 sky130_fd_sc_hd__nand2_1 _4384_ (.A(_3459_),
    .B(_0154_),
    .Y(_0158_));
 sky130_fd_sc_hd__o211ai_4 _4385_ (.A1(_0123_),
    .A2(_0126_),
    .B1(_0157_),
    .C1(_0158_),
    .Y(_0159_));
 sky130_fd_sc_hd__nand4_2 _4386_ (.A(net325),
    .B(net314),
    .C(net166),
    .D(net161),
    .Y(_0160_));
 sky130_fd_sc_hd__a21bo_1 _4387_ (.A1(_0160_),
    .A2(_3452_),
    .B1_N(_3453_),
    .X(_0161_));
 sky130_fd_sc_hd__nand4_2 _4388_ (.A(_3452_),
    .B(net173),
    .C(net302),
    .D(_0160_),
    .Y(_0162_));
 sky130_fd_sc_hd__nand2_1 _4389_ (.A(_0161_),
    .B(_0162_),
    .Y(_0163_));
 sky130_fd_sc_hd__nand2_4 _4390_ (.A(net337),
    .B(net166),
    .Y(_0164_));
 sky130_fd_sc_hd__nand2_1 _4391_ (.A(net173),
    .B(net314),
    .Y(_0165_));
 sky130_fd_sc_hd__a22oi_1 _4392_ (.A1(net327),
    .A2(net166),
    .B1(net161),
    .B2(net337),
    .Y(_0166_));
 sky130_fd_sc_hd__o22a_1 _4393_ (.A1(_3450_),
    .A2(_0164_),
    .B1(_0165_),
    .B2(_0166_),
    .X(_0167_));
 sky130_fd_sc_hd__o2bb2ai_2 _4394_ (.A1_N(_0156_),
    .A2_N(_0159_),
    .B1(_0163_),
    .B2(_0167_),
    .Y(_0168_));
 sky130_fd_sc_hd__nand4_1 _4395_ (.A(net337),
    .B(net325),
    .C(net166),
    .D(net161),
    .Y(_0169_));
 sky130_fd_sc_hd__o21ai_1 _4396_ (.A1(_0165_),
    .A2(_0166_),
    .B1(_0169_),
    .Y(_0170_));
 sky130_fd_sc_hd__and3_2 _4397_ (.A(_0161_),
    .B(_0162_),
    .C(_0170_),
    .X(_0171_));
 sky130_fd_sc_hd__nand3_2 _4398_ (.A(_0159_),
    .B(_0171_),
    .C(_0156_),
    .Y(_0172_));
 sky130_fd_sc_hd__nand3_1 _4399_ (.A(_0153_),
    .B(_0168_),
    .C(_0172_),
    .Y(_0173_));
 sky130_fd_sc_hd__nand3_1 _4400_ (.A(_3500_),
    .B(_3486_),
    .C(_3501_),
    .Y(_0174_));
 sky130_fd_sc_hd__a21o_1 _4401_ (.A1(_3500_),
    .A2(_3486_),
    .B1(_3501_),
    .X(_0175_));
 sky130_fd_sc_hd__nand4_2 _4402_ (.A(_0150_),
    .B(_0173_),
    .C(_0174_),
    .D(_0175_),
    .Y(_0176_));
 sky130_fd_sc_hd__nand2_1 _4403_ (.A(_3500_),
    .B(_3486_),
    .Y(_0177_));
 sky130_fd_sc_hd__nand2_1 _4404_ (.A(_3501_),
    .B(_0177_),
    .Y(_0178_));
 sky130_fd_sc_hd__nand2_1 _4405_ (.A(_0150_),
    .B(_0173_),
    .Y(_0179_));
 sky130_fd_sc_hd__nand4_1 _4406_ (.A(_3465_),
    .B(_3500_),
    .C(_3486_),
    .D(_3490_),
    .Y(_0180_));
 sky130_fd_sc_hd__nand3_1 _4407_ (.A(_0178_),
    .B(_0179_),
    .C(_0180_),
    .Y(_0181_));
 sky130_fd_sc_hd__a21boi_2 _4408_ (.A1(_0159_),
    .A2(_0171_),
    .B1_N(_0156_),
    .Y(_0182_));
 sky130_fd_sc_hd__nand2_1 _4409_ (.A(_0181_),
    .B(_0182_),
    .Y(_0183_));
 sky130_fd_sc_hd__nand2_1 _4410_ (.A(_0176_),
    .B(_0183_),
    .Y(_0184_));
 sky130_fd_sc_hd__a21oi_1 _4411_ (.A1(_0121_),
    .A2(_0122_),
    .B1(_0184_),
    .Y(_0185_));
 sky130_fd_sc_hd__a21oi_1 _4412_ (.A1(_3493_),
    .A2(_3503_),
    .B1(_3466_),
    .Y(_0186_));
 sky130_fd_sc_hd__nand2_1 _4413_ (.A(_0122_),
    .B(_0184_),
    .Y(_0187_));
 sky130_fd_sc_hd__a21o_1 _4414_ (.A1(_0176_),
    .A2(_0181_),
    .B1(_0182_),
    .X(_0188_));
 sky130_fd_sc_hd__nand3_1 _4415_ (.A(_0176_),
    .B(_0181_),
    .C(_0182_),
    .Y(_0189_));
 sky130_fd_sc_hd__a21oi_1 _4416_ (.A1(_0156_),
    .A2(_0159_),
    .B1(_0171_),
    .Y(_0190_));
 sky130_fd_sc_hd__inv_2 _4417_ (.A(_0172_),
    .Y(_0191_));
 sky130_fd_sc_hd__o2bb2ai_1 _4418_ (.A1_N(_0153_),
    .A2_N(_0150_),
    .B1(_0190_),
    .B2(_0191_),
    .Y(_0192_));
 sky130_fd_sc_hd__nand4_1 _4419_ (.A(_0153_),
    .B(_0150_),
    .C(_0168_),
    .D(_0172_),
    .Y(_0193_));
 sky130_fd_sc_hd__a21oi_2 _4420_ (.A1(_0144_),
    .A2(_0137_),
    .B1(_0141_),
    .Y(_0194_));
 sky130_fd_sc_hd__nand2_1 _4421_ (.A(net371),
    .B(net141),
    .Y(_0195_));
 sky130_fd_sc_hd__nand2_1 _4422_ (.A(_3442_),
    .B(_0195_),
    .Y(_0196_));
 sky130_fd_sc_hd__o21ai_1 _4423_ (.A1(_2555_),
    .A2(_0133_),
    .B1(_0196_),
    .Y(_0197_));
 sky130_fd_sc_hd__nor2_1 _4424_ (.A(_1825_),
    .B(_3049_),
    .Y(_0198_));
 sky130_fd_sc_hd__nand2_1 _4425_ (.A(_0197_),
    .B(_0198_),
    .Y(_0199_));
 sky130_fd_sc_hd__nand4_2 _4426_ (.A(net382),
    .B(net376),
    .C(net148),
    .D(net141),
    .Y(_0200_));
 sky130_fd_sc_hd__nand2_1 _4427_ (.A(net364),
    .B(net154),
    .Y(_0201_));
 sky130_fd_sc_hd__a22oi_1 _4428_ (.A1(net376),
    .A2(net148),
    .B1(net141),
    .B2(net382),
    .Y(_0202_));
 sky130_fd_sc_hd__a21o_1 _4429_ (.A1(_0200_),
    .A2(_0201_),
    .B1(_0202_),
    .X(_0203_));
 sky130_fd_sc_hd__o221ai_2 _4430_ (.A1(_2965_),
    .A2(_3049_),
    .B1(_2555_),
    .B2(_0133_),
    .C1(_0196_),
    .Y(_0204_));
 sky130_fd_sc_hd__nand3_2 _4431_ (.A(_0199_),
    .B(_0203_),
    .C(_0204_),
    .Y(_0205_));
 sky130_fd_sc_hd__a41o_1 _4432_ (.A1(net371),
    .A2(net359),
    .A3(net148),
    .A4(net141),
    .B1(_0134_),
    .X(_0206_));
 sky130_fd_sc_hd__a21oi_1 _4433_ (.A1(_0200_),
    .A2(_0201_),
    .B1(_0202_),
    .Y(_0207_));
 sky130_fd_sc_hd__nand4_1 _4434_ (.A(net371),
    .B(net359),
    .C(net148),
    .D(net141),
    .Y(_0208_));
 sky130_fd_sc_hd__o2bb2ai_2 _4435_ (.A1_N(_0208_),
    .A2_N(_0196_),
    .B1(_2965_),
    .B2(_3049_),
    .Y(_0209_));
 sky130_fd_sc_hd__o211ai_4 _4436_ (.A1(_0135_),
    .A2(_0206_),
    .B1(_0207_),
    .C1(_0209_),
    .Y(_0210_));
 sky130_fd_sc_hd__a22oi_2 _4437_ (.A1(net384),
    .A2(net135),
    .B1(net127),
    .B2(net394),
    .Y(_0211_));
 sky130_fd_sc_hd__nor2_2 _4438_ (.A(_0125_),
    .B(_0211_),
    .Y(_0212_));
 sky130_fd_sc_hd__and3_1 _4439_ (.A(_0205_),
    .B(_0210_),
    .C(_0212_),
    .X(_0213_));
 sky130_fd_sc_hd__nand2_2 _4440_ (.A(_0145_),
    .B(_0213_),
    .Y(_0214_));
 sky130_fd_sc_hd__a21o_1 _4441_ (.A1(_0160_),
    .A2(_3452_),
    .B1(_3453_),
    .X(_0215_));
 sky130_fd_sc_hd__o211ai_1 _4442_ (.A1(_3022_),
    .A2(_3313_),
    .B1(_0160_),
    .C1(_3452_),
    .Y(_0216_));
 sky130_fd_sc_hd__nand3_1 _4443_ (.A(_0215_),
    .B(_0216_),
    .C(_0167_),
    .Y(_0217_));
 sky130_fd_sc_hd__nand3_2 _4444_ (.A(_0161_),
    .B(_0162_),
    .C(_0170_),
    .Y(_0218_));
 sky130_fd_sc_hd__nand3b_2 _4445_ (.A_N(_0210_),
    .B(_0217_),
    .C(_0218_),
    .Y(_0219_));
 sky130_fd_sc_hd__o21ai_1 _4446_ (.A1(_0135_),
    .A2(_0206_),
    .B1(_0209_),
    .Y(_0220_));
 sky130_fd_sc_hd__o2bb2ai_2 _4447_ (.A1_N(_0218_),
    .A2_N(_0217_),
    .B1(_0220_),
    .B2(_0203_),
    .Y(_0221_));
 sky130_fd_sc_hd__nand2_1 _4448_ (.A(_0219_),
    .B(_0221_),
    .Y(_0222_));
 sky130_fd_sc_hd__nand2_1 _4449_ (.A(net325),
    .B(net166),
    .Y(_0223_));
 sky130_fd_sc_hd__nand2_2 _4450_ (.A(net338),
    .B(net161),
    .Y(_0224_));
 sky130_fd_sc_hd__nand2_2 _4451_ (.A(_0223_),
    .B(_0224_),
    .Y(_0225_));
 sky130_fd_sc_hd__and2_1 _4452_ (.A(net173),
    .B(net314),
    .X(_0226_));
 sky130_fd_sc_hd__a21o_1 _4453_ (.A1(_0225_),
    .A2(_0169_),
    .B1(_0226_),
    .X(_0227_));
 sky130_fd_sc_hd__o2111ai_4 _4454_ (.A1(_3450_),
    .A2(_0164_),
    .B1(net173),
    .C1(net315),
    .D1(_0225_),
    .Y(_0228_));
 sky130_fd_sc_hd__nand2_4 _4455_ (.A(net351),
    .B(net159),
    .Y(_0229_));
 sky130_fd_sc_hd__nand4_2 _4456_ (.A(net351),
    .B(net337),
    .C(net166),
    .D(net160),
    .Y(_0230_));
 sky130_fd_sc_hd__nand2_1 _4457_ (.A(net172),
    .B(net325),
    .Y(_0231_));
 sky130_fd_sc_hd__a22oi_4 _4458_ (.A1(_0164_),
    .A2(_0229_),
    .B1(_0230_),
    .B2(_0231_),
    .Y(_0232_));
 sky130_fd_sc_hd__nand3_2 _4459_ (.A(_0227_),
    .B(_0228_),
    .C(_0232_),
    .Y(_0233_));
 sky130_fd_sc_hd__nand2_1 _4460_ (.A(_0222_),
    .B(_0233_),
    .Y(_0234_));
 sky130_fd_sc_hd__nand3b_2 _4461_ (.A_N(_0233_),
    .B(_0221_),
    .C(_0219_),
    .Y(_0235_));
 sky130_fd_sc_hd__nand2_1 _4462_ (.A(_0234_),
    .B(_0235_),
    .Y(_0236_));
 sky130_fd_sc_hd__and2_1 _4463_ (.A(_0205_),
    .B(_0210_),
    .X(_0237_));
 sky130_fd_sc_hd__a21o_1 _4464_ (.A1(_0143_),
    .A2(_0131_),
    .B1(_0136_),
    .X(_0238_));
 sky130_fd_sc_hd__nand3_1 _4465_ (.A(_0131_),
    .B(_0136_),
    .C(_0143_),
    .Y(_0239_));
 sky130_fd_sc_hd__nand3b_2 _4466_ (.A_N(_0141_),
    .B(_0238_),
    .C(_0239_),
    .Y(_0240_));
 sky130_fd_sc_hd__a22oi_4 _4467_ (.A1(_0212_),
    .A2(_0237_),
    .B1(_0240_),
    .B2(_0145_),
    .Y(_0241_));
 sky130_fd_sc_hd__o22ai_1 _4468_ (.A1(_0194_),
    .A2(_0214_),
    .B1(_0236_),
    .B2(_0241_),
    .Y(_0242_));
 sky130_fd_sc_hd__nand3_1 _4469_ (.A(_0192_),
    .B(_0193_),
    .C(_0242_),
    .Y(_0243_));
 sky130_fd_sc_hd__inv_2 _4470_ (.A(_0219_),
    .Y(_0244_));
 sky130_fd_sc_hd__a41o_1 _4471_ (.A1(_0221_),
    .A2(_0232_),
    .A3(_0227_),
    .A4(_0228_),
    .B1(_0244_),
    .X(_0245_));
 sky130_fd_sc_hd__inv_2 _4472_ (.A(_0245_),
    .Y(_0246_));
 sky130_fd_sc_hd__nand3_2 _4473_ (.A(_0205_),
    .B(_0210_),
    .C(_0212_),
    .Y(_0247_));
 sky130_fd_sc_hd__a31oi_1 _4474_ (.A1(_0137_),
    .A2(_0141_),
    .A3(_0144_),
    .B1(_0247_),
    .Y(_0248_));
 sky130_fd_sc_hd__a22oi_1 _4475_ (.A1(_0234_),
    .A2(_0235_),
    .B1(_0240_),
    .B2(_0248_),
    .Y(_0249_));
 sky130_fd_sc_hd__nand2_1 _4476_ (.A(_0168_),
    .B(_0172_),
    .Y(_0250_));
 sky130_fd_sc_hd__nand3_1 _4477_ (.A(_0153_),
    .B(_0150_),
    .C(_0250_),
    .Y(_0251_));
 sky130_fd_sc_hd__a21oi_1 _4478_ (.A1(_0156_),
    .A2(_0159_),
    .B1(_0218_),
    .Y(_0252_));
 sky130_fd_sc_hd__and3_1 _4479_ (.A(_0218_),
    .B(_0156_),
    .C(_0159_),
    .X(_0253_));
 sky130_fd_sc_hd__o2bb2ai_1 _4480_ (.A1_N(_0153_),
    .A2_N(_0150_),
    .B1(_0252_),
    .B2(_0253_),
    .Y(_0254_));
 sky130_fd_sc_hd__o211ai_2 _4481_ (.A1(_0241_),
    .A2(_0249_),
    .B1(_0251_),
    .C1(_0254_),
    .Y(_0255_));
 sky130_fd_sc_hd__a21bo_1 _4482_ (.A1(_0243_),
    .A2(_0246_),
    .B1_N(_0255_),
    .X(_0256_));
 sky130_fd_sc_hd__nand3_1 _4483_ (.A(_0188_),
    .B(_0189_),
    .C(_0256_),
    .Y(_0257_));
 sky130_fd_sc_hd__o21a_1 _4484_ (.A1(_0186_),
    .A2(_0187_),
    .B1(_0257_),
    .X(_0258_));
 sky130_fd_sc_hd__a21o_1 _4485_ (.A1(_0121_),
    .A2(_0122_),
    .B1(_0184_),
    .X(_0259_));
 sky130_fd_sc_hd__nand2_1 _4486_ (.A(_0176_),
    .B(_0181_),
    .Y(_0260_));
 sky130_fd_sc_hd__and4_1 _4487_ (.A(_0221_),
    .B(_0232_),
    .C(_0227_),
    .D(_0228_),
    .X(_0261_));
 sky130_fd_sc_hd__o21ai_1 _4488_ (.A1(_0244_),
    .A2(_0261_),
    .B1(_0255_),
    .Y(_0262_));
 sky130_fd_sc_hd__a22oi_1 _4489_ (.A1(_0243_),
    .A2(_0262_),
    .B1(_0260_),
    .B2(_0182_),
    .Y(_0263_));
 sky130_fd_sc_hd__o21ai_1 _4490_ (.A1(_0182_),
    .A2(_0260_),
    .B1(_0263_),
    .Y(_0264_));
 sky130_fd_sc_hd__nand2_1 _4491_ (.A(_0259_),
    .B(_0264_),
    .Y(_0265_));
 sky130_fd_sc_hd__nor2_1 _4492_ (.A(_0194_),
    .B(_0214_),
    .Y(_0266_));
 sky130_fd_sc_hd__o21ai_1 _4493_ (.A1(_0241_),
    .A2(_0266_),
    .B1(_0236_),
    .Y(_0267_));
 sky130_fd_sc_hd__nand2_1 _4494_ (.A(_0205_),
    .B(_0210_),
    .Y(_0268_));
 sky130_fd_sc_hd__inv_2 _4495_ (.A(_0212_),
    .Y(_0269_));
 sky130_fd_sc_hd__o2bb2ai_2 _4496_ (.A1_N(_0145_),
    .A2_N(_0240_),
    .B1(_0268_),
    .B2(_0269_),
    .Y(_0270_));
 sky130_fd_sc_hd__o2111ai_4 _4497_ (.A1(_0194_),
    .A2(_0214_),
    .B1(_0234_),
    .C1(_0235_),
    .D1(_0270_),
    .Y(_0271_));
 sky130_fd_sc_hd__nand2_1 _4498_ (.A(net376),
    .B(net148),
    .Y(_0272_));
 sky130_fd_sc_hd__nand2_1 _4499_ (.A(net385),
    .B(net141),
    .Y(_0273_));
 sky130_fd_sc_hd__nand2_1 _4500_ (.A(_0272_),
    .B(_0273_),
    .Y(_0274_));
 sky130_fd_sc_hd__o2bb2ai_2 _4501_ (.A1_N(_0200_),
    .A2_N(_0274_),
    .B1(_1727_),
    .B2(_3049_),
    .Y(_0275_));
 sky130_fd_sc_hd__nand4_2 _4502_ (.A(_0274_),
    .B(net154),
    .C(net364),
    .D(_0200_),
    .Y(_0276_));
 sky130_fd_sc_hd__nand2_1 _4503_ (.A(net375),
    .B(net154),
    .Y(_0277_));
 sky130_fd_sc_hd__a22oi_1 _4504_ (.A1(net386),
    .A2(net149),
    .B1(net142),
    .B2(net396),
    .Y(_0278_));
 sky130_fd_sc_hd__nand4_4 _4505_ (.A(net396),
    .B(net386),
    .C(net149),
    .D(net142),
    .Y(_0279_));
 sky130_fd_sc_hd__o21ai_1 _4506_ (.A1(_0277_),
    .A2(_0278_),
    .B1(_0279_),
    .Y(_0280_));
 sky130_fd_sc_hd__nand3_1 _4507_ (.A(_0275_),
    .B(_0276_),
    .C(_0280_),
    .Y(_0281_));
 sky130_fd_sc_hd__a22o_1 _4508_ (.A1(_0164_),
    .A2(_0229_),
    .B1(_0230_),
    .B2(_0231_),
    .X(_0282_));
 sky130_fd_sc_hd__o221ai_1 _4509_ (.A1(_3313_),
    .A2(_2794_),
    .B1(_3450_),
    .B2(_0164_),
    .C1(_0225_),
    .Y(_0283_));
 sky130_fd_sc_hd__nand2_1 _4510_ (.A(_0225_),
    .B(_0169_),
    .Y(_0284_));
 sky130_fd_sc_hd__nand2_1 _4511_ (.A(_0284_),
    .B(_0226_),
    .Y(_0285_));
 sky130_fd_sc_hd__nand3_1 _4512_ (.A(_0282_),
    .B(_0283_),
    .C(_0285_),
    .Y(_0286_));
 sky130_fd_sc_hd__nand3b_1 _4513_ (.A_N(_0281_),
    .B(_0286_),
    .C(_0233_),
    .Y(_0287_));
 sky130_fd_sc_hd__nand2_1 _4514_ (.A(_0275_),
    .B(_0276_),
    .Y(_0288_));
 sky130_fd_sc_hd__o31a_1 _4515_ (.A1(_2218_),
    .A2(_1445_),
    .A3(_0278_),
    .B1(_0279_),
    .X(_0289_));
 sky130_fd_sc_hd__o2bb2ai_1 _4516_ (.A1_N(_0233_),
    .A2_N(_0286_),
    .B1(_0288_),
    .B2(_0289_),
    .Y(_0290_));
 sky130_fd_sc_hd__clkbuf_2 _4517_ (.A(_0290_),
    .X(_0291_));
 sky130_fd_sc_hd__nand2_2 _4518_ (.A(net363),
    .B(net168),
    .Y(_0292_));
 sky130_fd_sc_hd__nand2_1 _4519_ (.A(net171),
    .B(net337),
    .Y(_0293_));
 sky130_fd_sc_hd__a22oi_2 _4520_ (.A1(net351),
    .A2(net167),
    .B1(net159),
    .B2(net363),
    .Y(_0294_));
 sky130_fd_sc_hd__o22a_1 _4521_ (.A1(_0229_),
    .A2(_0292_),
    .B1(_0293_),
    .B2(_0294_),
    .X(_0295_));
 sky130_fd_sc_hd__nand2_2 _4522_ (.A(_0164_),
    .B(_0229_),
    .Y(_0296_));
 sky130_fd_sc_hd__a22o_2 _4523_ (.A1(net172),
    .A2(net325),
    .B1(_0296_),
    .B2(_0230_),
    .X(_0297_));
 sky130_fd_sc_hd__nand2_2 _4524_ (.A(net351),
    .B(net168),
    .Y(_0298_));
 sky130_fd_sc_hd__o2111ai_4 _4525_ (.A1(_0224_),
    .A2(_0298_),
    .B1(net173),
    .C1(net325),
    .D1(_0296_),
    .Y(_0299_));
 sky130_fd_sc_hd__nand2_1 _4526_ (.A(_0297_),
    .B(_0299_),
    .Y(_0300_));
 sky130_fd_sc_hd__o2bb2ai_1 _4527_ (.A1_N(_0287_),
    .A2_N(_0291_),
    .B1(_0295_),
    .B2(_0300_),
    .Y(_0301_));
 sky130_fd_sc_hd__nand4_4 _4528_ (.A(net363),
    .B(net351),
    .C(net167),
    .D(net159),
    .Y(_0302_));
 sky130_fd_sc_hd__o21ai_4 _4529_ (.A1(_0293_),
    .A2(_0294_),
    .B1(_0302_),
    .Y(_0303_));
 sky130_fd_sc_hd__nand3_4 _4530_ (.A(_0297_),
    .B(_0299_),
    .C(_0303_),
    .Y(_0304_));
 sky130_fd_sc_hd__clkbuf_2 _4531_ (.A(_0287_),
    .X(_0305_));
 sky130_fd_sc_hd__nand3b_1 _4532_ (.A_N(_0304_),
    .B(_0291_),
    .C(_0305_),
    .Y(_0306_));
 sky130_fd_sc_hd__nand2_1 _4533_ (.A(_0301_),
    .B(_0306_),
    .Y(_0307_));
 sky130_fd_sc_hd__a21o_2 _4534_ (.A1(_0275_),
    .A2(_0276_),
    .B1(_0280_),
    .X(_0308_));
 sky130_fd_sc_hd__and3_1 _4535_ (.A(_0281_),
    .B(net134),
    .C(net394),
    .X(_0309_));
 sky130_fd_sc_hd__a21oi_1 _4536_ (.A1(_0205_),
    .A2(_0210_),
    .B1(_0212_),
    .Y(_0310_));
 sky130_fd_sc_hd__o2bb2ai_2 _4537_ (.A1_N(_0308_),
    .A2_N(_0309_),
    .B1(_0310_),
    .B2(_0213_),
    .Y(_0311_));
 sky130_fd_sc_hd__inv_2 _4538_ (.A(_0311_),
    .Y(_0312_));
 sky130_fd_sc_hd__o21ai_2 _4539_ (.A1(_0125_),
    .A2(_0211_),
    .B1(_0268_),
    .Y(_0313_));
 sky130_fd_sc_hd__nand4_4 _4540_ (.A(_0309_),
    .B(_0313_),
    .C(_0247_),
    .D(_0308_),
    .Y(_0314_));
 sky130_fd_sc_hd__o21ai_1 _4541_ (.A1(_0307_),
    .A2(_0312_),
    .B1(_0314_),
    .Y(_0315_));
 sky130_fd_sc_hd__o21bai_1 _4542_ (.A1(_0241_),
    .A2(_0266_),
    .B1_N(_0236_),
    .Y(_0316_));
 sky130_fd_sc_hd__o211ai_1 _4543_ (.A1(_0194_),
    .A2(_0214_),
    .B1(_0236_),
    .C1(_0270_),
    .Y(_0317_));
 sky130_fd_sc_hd__a21o_1 _4544_ (.A1(_0305_),
    .A2(_0291_),
    .B1(_0304_),
    .X(_0318_));
 sky130_fd_sc_hd__o211ai_2 _4545_ (.A1(_0295_),
    .A2(_0300_),
    .B1(_0305_),
    .C1(_0291_),
    .Y(_0319_));
 sky130_fd_sc_hd__a31o_1 _4546_ (.A1(_0314_),
    .A2(_0318_),
    .A3(_0319_),
    .B1(_0312_),
    .X(_0320_));
 sky130_fd_sc_hd__nand3_2 _4547_ (.A(_0316_),
    .B(_0317_),
    .C(_0320_),
    .Y(_0321_));
 sky130_fd_sc_hd__inv_2 _4548_ (.A(_0305_),
    .Y(_0322_));
 sky130_fd_sc_hd__a41o_1 _4549_ (.A1(_0291_),
    .A2(_0303_),
    .A3(_0297_),
    .A4(_0299_),
    .B1(_0322_),
    .X(_0323_));
 sky130_fd_sc_hd__a32o_1 _4550_ (.A1(_0267_),
    .A2(_0271_),
    .A3(_0315_),
    .B1(_0321_),
    .B2(_0323_),
    .X(_0324_));
 sky130_fd_sc_hd__o2bb2ai_1 _4551_ (.A1_N(_0243_),
    .A2_N(_0255_),
    .B1(_0261_),
    .B2(_0244_),
    .Y(_0325_));
 sky130_fd_sc_hd__nand3_1 _4552_ (.A(_0243_),
    .B(_0255_),
    .C(_0246_),
    .Y(_0326_));
 sky130_fd_sc_hd__nand2_1 _4553_ (.A(_0325_),
    .B(_0326_),
    .Y(_0327_));
 sky130_fd_sc_hd__o2bb2a_1 _4554_ (.A1_N(_0233_),
    .A2_N(_0286_),
    .B1(_0288_),
    .B2(_0289_),
    .X(_0328_));
 sky130_fd_sc_hd__nand3_2 _4555_ (.A(_0267_),
    .B(_0271_),
    .C(_0315_),
    .Y(_0329_));
 sky130_fd_sc_hd__o2111ai_1 _4556_ (.A1(_0304_),
    .A2(_0328_),
    .B1(_0305_),
    .C1(_0321_),
    .D1(_0329_),
    .Y(_0330_));
 sky130_fd_sc_hd__and4_1 _4557_ (.A(_0291_),
    .B(_0303_),
    .C(_0297_),
    .D(_0299_),
    .X(_0331_));
 sky130_fd_sc_hd__o2bb2ai_1 _4558_ (.A1_N(_0329_),
    .A2_N(_0321_),
    .B1(_0331_),
    .B2(_0322_),
    .Y(_0332_));
 sky130_fd_sc_hd__o221ai_2 _4559_ (.A1(_3313_),
    .A2(_2886_),
    .B1(_0224_),
    .B2(_0298_),
    .C1(_0296_),
    .Y(_0333_));
 sky130_fd_sc_hd__o2bb2ai_1 _4560_ (.A1_N(_0164_),
    .A2_N(_0229_),
    .B1(_0298_),
    .B2(_0224_),
    .Y(_0334_));
 sky130_fd_sc_hd__nand3_1 _4561_ (.A(_0334_),
    .B(net325),
    .C(net172),
    .Y(_0335_));
 sky130_fd_sc_hd__nand3_2 _4562_ (.A(_0295_),
    .B(_0333_),
    .C(_0335_),
    .Y(_0336_));
 sky130_fd_sc_hd__nand2_1 _4563_ (.A(net386),
    .B(net149),
    .Y(_0337_));
 sky130_fd_sc_hd__nand2_1 _4564_ (.A(net396),
    .B(net142),
    .Y(_0338_));
 sky130_fd_sc_hd__a21oi_1 _4565_ (.A1(_0337_),
    .A2(_0338_),
    .B1(_0277_),
    .Y(_0339_));
 sky130_fd_sc_hd__nand4_1 _4566_ (.A(net396),
    .B(net386),
    .C(net153),
    .D(net148),
    .Y(_0340_));
 sky130_fd_sc_hd__nand2_1 _4567_ (.A(_0337_),
    .B(_0338_),
    .Y(_0341_));
 sky130_fd_sc_hd__a22oi_2 _4568_ (.A1(net375),
    .A2(net153),
    .B1(_0341_),
    .B2(_0279_),
    .Y(_0342_));
 sky130_fd_sc_hd__a211oi_2 _4569_ (.A1(_0279_),
    .A2(_0339_),
    .B1(_0340_),
    .C1(_0342_),
    .Y(_0343_));
 sky130_fd_sc_hd__a21oi_2 _4570_ (.A1(_0304_),
    .A2(_0336_),
    .B1(_0343_),
    .Y(_0344_));
 sky130_fd_sc_hd__o2bb2a_1 _4571_ (.A1_N(_0296_),
    .A2_N(_0230_),
    .B1(_3178_),
    .B2(_1793_),
    .X(_0345_));
 sky130_fd_sc_hd__o21ai_1 _4572_ (.A1(_0231_),
    .A2(_0334_),
    .B1(_0303_),
    .Y(_0346_));
 sky130_fd_sc_hd__o211ai_2 _4573_ (.A1(_0345_),
    .A2(_0346_),
    .B1(_0336_),
    .C1(_0343_),
    .Y(_0347_));
 sky130_fd_sc_hd__nand2_1 _4574_ (.A(net172),
    .B(net352),
    .Y(_0348_));
 sky130_fd_sc_hd__a22oi_4 _4575_ (.A1(net364),
    .A2(net168),
    .B1(net160),
    .B2(net375),
    .Y(_0349_));
 sky130_fd_sc_hd__nand4_4 _4576_ (.A(net376),
    .B(net364),
    .C(net167),
    .D(net159),
    .Y(_0350_));
 sky130_fd_sc_hd__o21ai_1 _4577_ (.A1(_0348_),
    .A2(_0349_),
    .B1(_0350_),
    .Y(_0351_));
 sky130_fd_sc_hd__nand2_1 _4578_ (.A(net363),
    .B(net161),
    .Y(_0352_));
 sky130_fd_sc_hd__nand2_2 _4579_ (.A(_0298_),
    .B(_0352_),
    .Y(_0353_));
 sky130_fd_sc_hd__a22oi_4 _4580_ (.A1(net171),
    .A2(net337),
    .B1(_0353_),
    .B2(_0302_),
    .Y(_0354_));
 sky130_fd_sc_hd__and2_1 _4581_ (.A(net171),
    .B(net338),
    .X(_0355_));
 sky130_fd_sc_hd__o211a_1 _4582_ (.A1(_0229_),
    .A2(_0292_),
    .B1(_0355_),
    .C1(_0353_),
    .X(_0356_));
 sky130_fd_sc_hd__nor2_1 _4583_ (.A(_0354_),
    .B(_0356_),
    .Y(_0357_));
 sky130_fd_sc_hd__nand4b_1 _4584_ (.A_N(_0344_),
    .B(_0347_),
    .C(_0351_),
    .D(_0357_),
    .Y(_0358_));
 sky130_fd_sc_hd__o2111ai_2 _4585_ (.A1(_0229_),
    .A2(_0292_),
    .B1(net173),
    .C1(net337),
    .D1(_0353_),
    .Y(_0359_));
 sky130_fd_sc_hd__nand2_1 _4586_ (.A(_0359_),
    .B(_0351_),
    .Y(_0360_));
 sky130_fd_sc_hd__o211a_1 _4587_ (.A1(_0345_),
    .A2(_0346_),
    .B1(_0336_),
    .C1(_0343_),
    .X(_0361_));
 sky130_fd_sc_hd__o22ai_2 _4588_ (.A1(_0354_),
    .A2(_0360_),
    .B1(_0344_),
    .B2(_0361_),
    .Y(_0362_));
 sky130_fd_sc_hd__a22oi_1 _4589_ (.A1(net394),
    .A2(net134),
    .B1(_0308_),
    .B2(_0281_),
    .Y(_0363_));
 sky130_fd_sc_hd__a21oi_1 _4590_ (.A1(_0308_),
    .A2(_0309_),
    .B1(_0363_),
    .Y(_0364_));
 sky130_fd_sc_hd__nand3_2 _4591_ (.A(_0358_),
    .B(_0362_),
    .C(_0364_),
    .Y(_0365_));
 sky130_fd_sc_hd__a21oi_1 _4592_ (.A1(_0305_),
    .A2(_0291_),
    .B1(_0304_),
    .Y(_0366_));
 sky130_fd_sc_hd__and3_1 _4593_ (.A(_0305_),
    .B(_0290_),
    .C(_0304_),
    .X(_0367_));
 sky130_fd_sc_hd__nand2_1 _4594_ (.A(_0311_),
    .B(_0314_),
    .Y(_0368_));
 sky130_fd_sc_hd__o21ai_1 _4595_ (.A1(_0366_),
    .A2(_0367_),
    .B1(_0368_),
    .Y(_0369_));
 sky130_fd_sc_hd__nand4_1 _4596_ (.A(_0311_),
    .B(_0314_),
    .C(_0318_),
    .D(_0319_),
    .Y(_0370_));
 sky130_fd_sc_hd__nand3_1 _4597_ (.A(_0365_),
    .B(_0369_),
    .C(_0370_),
    .Y(_0371_));
 sky130_fd_sc_hd__nand3b_1 _4598_ (.A_N(_0354_),
    .B(_0359_),
    .C(_0351_),
    .Y(_0372_));
 sky130_fd_sc_hd__o21ai_1 _4599_ (.A1(_0372_),
    .A2(_0344_),
    .B1(_0347_),
    .Y(_0373_));
 sky130_fd_sc_hd__nand2_1 _4600_ (.A(_0307_),
    .B(_0368_),
    .Y(_0374_));
 sky130_fd_sc_hd__nand4_1 _4601_ (.A(_0311_),
    .B(_0314_),
    .C(_0301_),
    .D(_0306_),
    .Y(_0375_));
 sky130_fd_sc_hd__nand3b_2 _4602_ (.A_N(_0365_),
    .B(_0374_),
    .C(_0375_),
    .Y(_0376_));
 sky130_fd_sc_hd__a21boi_1 _4603_ (.A1(_0371_),
    .A2(_0373_),
    .B1_N(_0376_),
    .Y(_0377_));
 sky130_fd_sc_hd__nand3_1 _4604_ (.A(_0330_),
    .B(_0332_),
    .C(_0377_),
    .Y(_0378_));
 sky130_fd_sc_hd__a21o_1 _4605_ (.A1(_0358_),
    .A2(_0362_),
    .B1(_0364_),
    .X(_0379_));
 sky130_fd_sc_hd__nand2_1 _4606_ (.A(net375),
    .B(net167),
    .Y(_0380_));
 sky130_fd_sc_hd__nand2_1 _4607_ (.A(net387),
    .B(net160),
    .Y(_0381_));
 sky130_fd_sc_hd__nand4_2 _4608_ (.A(net387),
    .B(net375),
    .C(net167),
    .D(net159),
    .Y(_0382_));
 sky130_fd_sc_hd__nand2_1 _4609_ (.A(net171),
    .B(net363),
    .Y(_0383_));
 sky130_fd_sc_hd__a22oi_2 _4610_ (.A1(_0380_),
    .A2(_0381_),
    .B1(_0382_),
    .B2(_0383_),
    .Y(_0384_));
 sky130_fd_sc_hd__buf_4 _4611_ (.A(_1825_),
    .X(_0385_));
 sky130_fd_sc_hd__nand2_1 _4612_ (.A(net375),
    .B(net161),
    .Y(_0386_));
 sky130_fd_sc_hd__nand3_1 _4613_ (.A(_0386_),
    .B(net168),
    .C(net363),
    .Y(_0387_));
 sky130_fd_sc_hd__nand3_1 _4614_ (.A(_0292_),
    .B(net161),
    .C(net375),
    .Y(_0388_));
 sky130_fd_sc_hd__o211ai_2 _4615_ (.A1(_3313_),
    .A2(_0385_),
    .B1(_0387_),
    .C1(_0388_),
    .Y(_0389_));
 sky130_fd_sc_hd__nand2_1 _4616_ (.A(_0292_),
    .B(_0386_),
    .Y(_0390_));
 sky130_fd_sc_hd__nand4_2 _4617_ (.A(_0390_),
    .B(_0350_),
    .C(net172),
    .D(net351),
    .Y(_0391_));
 sky130_fd_sc_hd__o221ai_4 _4618_ (.A1(_0349_),
    .A2(_0348_),
    .B1(_0354_),
    .B2(_0356_),
    .C1(_0350_),
    .Y(_0392_));
 sky130_fd_sc_hd__a32o_1 _4619_ (.A1(_0384_),
    .A2(_0389_),
    .A3(_0391_),
    .B1(_0392_),
    .B2(_0372_),
    .X(_0393_));
 sky130_fd_sc_hd__and3_1 _4620_ (.A(_0389_),
    .B(_0391_),
    .C(_0384_),
    .X(_0394_));
 sky130_fd_sc_hd__nor2_2 _4621_ (.A(_3125_),
    .B(_3050_),
    .Y(_0395_));
 sky130_fd_sc_hd__a21oi_1 _4622_ (.A1(_0279_),
    .A2(_0339_),
    .B1(_0342_),
    .Y(_0396_));
 sky130_fd_sc_hd__a31oi_1 _4623_ (.A1(net386),
    .A2(net149),
    .A3(_0395_),
    .B1(_0396_),
    .Y(_0397_));
 sky130_fd_sc_hd__nor2_1 _4624_ (.A(_0343_),
    .B(_0397_),
    .Y(_0398_));
 sky130_fd_sc_hd__a31o_1 _4625_ (.A1(_0372_),
    .A2(_0394_),
    .A3(_0392_),
    .B1(_0398_),
    .X(_0399_));
 sky130_fd_sc_hd__nand4_2 _4626_ (.A(_0365_),
    .B(_0379_),
    .C(_0393_),
    .D(_0399_),
    .Y(_0400_));
 sky130_fd_sc_hd__o211ai_2 _4627_ (.A1(_0354_),
    .A2(_0360_),
    .B1(_0394_),
    .C1(_0392_),
    .Y(_0401_));
 sky130_fd_sc_hd__nand2_1 _4628_ (.A(_0393_),
    .B(_0401_),
    .Y(_0402_));
 sky130_fd_sc_hd__a22oi_2 _4629_ (.A1(net386),
    .A2(net153),
    .B1(net149),
    .B2(net397),
    .Y(_0403_));
 sky130_fd_sc_hd__a31o_1 _4630_ (.A1(net386),
    .A2(net149),
    .A3(_0395_),
    .B1(_0403_),
    .X(_0404_));
 sky130_fd_sc_hd__nand3_1 _4631_ (.A(_0389_),
    .B(_0391_),
    .C(_0384_),
    .Y(_0405_));
 sky130_fd_sc_hd__a21o_1 _4632_ (.A1(_0389_),
    .A2(_0391_),
    .B1(_0384_),
    .X(_0406_));
 sky130_fd_sc_hd__nand2_1 _4633_ (.A(_0380_),
    .B(_0381_),
    .Y(_0407_));
 sky130_fd_sc_hd__nand4_2 _4634_ (.A(_0407_),
    .B(_0382_),
    .C(net171),
    .D(net363),
    .Y(_0408_));
 sky130_fd_sc_hd__nand2_1 _4635_ (.A(net172),
    .B(net375),
    .Y(_0409_));
 sky130_fd_sc_hd__a22oi_1 _4636_ (.A1(net387),
    .A2(net167),
    .B1(net159),
    .B2(net396),
    .Y(_0410_));
 sky130_fd_sc_hd__nand4_1 _4637_ (.A(net396),
    .B(net387),
    .C(net167),
    .D(net159),
    .Y(_0411_));
 sky130_fd_sc_hd__o21ai_2 _4638_ (.A1(_0409_),
    .A2(_0410_),
    .B1(_0411_),
    .Y(_0412_));
 sky130_fd_sc_hd__nand2_1 _4639_ (.A(_0408_),
    .B(_0412_),
    .Y(_0413_));
 sky130_fd_sc_hd__o2bb2a_1 _4640_ (.A1_N(_0407_),
    .A2_N(_0382_),
    .B1(_3178_),
    .B2(_3134_),
    .X(_0414_));
 sky130_fd_sc_hd__o2bb2a_1 _4641_ (.A1_N(_0405_),
    .A2_N(_0406_),
    .B1(_0413_),
    .B2(_0414_),
    .X(_0415_));
 sky130_fd_sc_hd__a22o_1 _4642_ (.A1(net171),
    .A2(net363),
    .B1(_0407_),
    .B2(_0382_),
    .X(_0416_));
 sky130_fd_sc_hd__and3_1 _4643_ (.A(_0416_),
    .B(_0408_),
    .C(_0412_),
    .X(_0417_));
 sky130_fd_sc_hd__nand3_1 _4644_ (.A(_0417_),
    .B(_0406_),
    .C(_0405_),
    .Y(_0418_));
 sky130_fd_sc_hd__o21ai_1 _4645_ (.A1(_0404_),
    .A2(_0415_),
    .B1(_0418_),
    .Y(_0419_));
 sky130_fd_sc_hd__a21oi_1 _4646_ (.A1(_0402_),
    .A2(_0398_),
    .B1(_0419_),
    .Y(_0420_));
 sky130_fd_sc_hd__or2_1 _4647_ (.A(_0398_),
    .B(_0402_),
    .X(_0421_));
 sky130_fd_sc_hd__a32o_1 _4648_ (.A1(_0412_),
    .A2(_0416_),
    .A3(_0408_),
    .B1(_0406_),
    .B2(_0405_),
    .X(_0422_));
 sky130_fd_sc_hd__nand2_1 _4649_ (.A(_0418_),
    .B(_0422_),
    .Y(_0423_));
 sky130_fd_sc_hd__nor2_1 _4650_ (.A(_3177_),
    .B(_3124_),
    .Y(_0057_));
 sky130_fd_sc_hd__and3_1 _4651_ (.A(net387),
    .B(net167),
    .C(_0057_),
    .X(_0424_));
 sky130_fd_sc_hd__clkbuf_2 _4652_ (.A(_0424_),
    .X(_0425_));
 sky130_fd_sc_hd__a22o_1 _4653_ (.A1(net387),
    .A2(net168),
    .B1(net159),
    .B2(net396),
    .X(_0426_));
 sky130_fd_sc_hd__and3_1 _4654_ (.A(_0411_),
    .B(net376),
    .C(net171),
    .X(_0427_));
 sky130_fd_sc_hd__a22oi_1 _4655_ (.A1(net171),
    .A2(net376),
    .B1(_0426_),
    .B2(_0411_),
    .Y(_0428_));
 sky130_fd_sc_hd__a21oi_2 _4656_ (.A1(_0426_),
    .A2(_0427_),
    .B1(_0428_),
    .Y(_0429_));
 sky130_fd_sc_hd__a21oi_1 _4657_ (.A1(_0416_),
    .A2(_0408_),
    .B1(_0412_),
    .Y(_0430_));
 sky130_fd_sc_hd__o2bb2ai_1 _4658_ (.A1_N(_0425_),
    .A2_N(_0429_),
    .B1(_0430_),
    .B2(_0417_),
    .Y(_0431_));
 sky130_fd_sc_hd__o211ai_1 _4659_ (.A1(_0414_),
    .A2(_0413_),
    .B1(_0425_),
    .C1(_0429_),
    .Y(_0432_));
 sky130_fd_sc_hd__o2bb2ai_1 _4660_ (.A1_N(_0395_),
    .A2_N(_0431_),
    .B1(_0432_),
    .B2(_0430_),
    .Y(_0433_));
 sky130_fd_sc_hd__o21a_1 _4661_ (.A1(_0404_),
    .A2(_0423_),
    .B1(_0433_),
    .X(_0434_));
 sky130_fd_sc_hd__nand2_1 _4662_ (.A(_0404_),
    .B(_0423_),
    .Y(_0435_));
 sky130_fd_sc_hd__nand2_1 _4663_ (.A(_0434_),
    .B(_0435_),
    .Y(_0436_));
 sky130_fd_sc_hd__nand3_1 _4664_ (.A(_0393_),
    .B(_0401_),
    .C(_0398_),
    .Y(_0437_));
 sky130_fd_sc_hd__a21o_1 _4665_ (.A1(_0393_),
    .A2(_0401_),
    .B1(_0398_),
    .X(_0438_));
 sky130_fd_sc_hd__nand3_1 _4666_ (.A(_0437_),
    .B(_0438_),
    .C(_0419_),
    .Y(_0439_));
 sky130_fd_sc_hd__a22oi_2 _4667_ (.A1(_0420_),
    .A2(_0421_),
    .B1(_0436_),
    .B2(_0439_),
    .Y(_0440_));
 sky130_fd_sc_hd__a22o_1 _4668_ (.A1(_0365_),
    .A2(_0379_),
    .B1(_0393_),
    .B2(_0399_),
    .X(_0441_));
 sky130_fd_sc_hd__nand2_1 _4669_ (.A(_0440_),
    .B(_0441_),
    .Y(_0442_));
 sky130_fd_sc_hd__nand3_1 _4670_ (.A(_0371_),
    .B(_0376_),
    .C(_0373_),
    .Y(_0443_));
 sky130_fd_sc_hd__o21a_1 _4671_ (.A1(_0354_),
    .A2(_0360_),
    .B1(_0347_),
    .X(_0444_));
 sky130_fd_sc_hd__o2bb2ai_1 _4672_ (.A1_N(_0371_),
    .A2_N(_0376_),
    .B1(_0444_),
    .B2(_0344_),
    .Y(_0445_));
 sky130_fd_sc_hd__nand2_1 _4673_ (.A(_0443_),
    .B(_0445_),
    .Y(_0446_));
 sky130_fd_sc_hd__a21oi_2 _4674_ (.A1(_0400_),
    .A2(_0442_),
    .B1(_0446_),
    .Y(_0447_));
 sky130_fd_sc_hd__nand2_2 _4675_ (.A(_0378_),
    .B(_0447_),
    .Y(_0448_));
 sky130_fd_sc_hd__a31oi_1 _4676_ (.A1(_0329_),
    .A2(_0321_),
    .A3(_0323_),
    .B1(_0377_),
    .Y(_0449_));
 sky130_fd_sc_hd__a21o_1 _4677_ (.A1(_0329_),
    .A2(_0321_),
    .B1(_0323_),
    .X(_0450_));
 sky130_fd_sc_hd__a22oi_2 _4678_ (.A1(_0449_),
    .A2(_0450_),
    .B1(_0327_),
    .B2(_0324_),
    .Y(_0451_));
 sky130_fd_sc_hd__a2bb2oi_4 _4679_ (.A1_N(_0324_),
    .A2_N(_0327_),
    .B1(_0448_),
    .B2(_0451_),
    .Y(_0452_));
 sky130_fd_sc_hd__o22ai_4 _4680_ (.A1(_0185_),
    .A2(_0258_),
    .B1(_0265_),
    .B2(_0452_),
    .Y(_0453_));
 sky130_fd_sc_hd__nand2_1 _4681_ (.A(_3506_),
    .B(_0119_),
    .Y(_0454_));
 sky130_fd_sc_hd__nand2_1 _4682_ (.A(_3533_),
    .B(_0106_),
    .Y(_0455_));
 sky130_fd_sc_hd__nand2_1 _4683_ (.A(_3528_),
    .B(_0455_),
    .Y(_0456_));
 sky130_fd_sc_hd__inv_2 _4684_ (.A(_3161_),
    .Y(_0457_));
 sky130_fd_sc_hd__o211ai_2 _4685_ (.A1(_3165_),
    .A2(_3164_),
    .B1(_3159_),
    .C1(_0457_),
    .Y(_0458_));
 sky130_fd_sc_hd__o21ai_1 _4686_ (.A1(_3165_),
    .A2(_3164_),
    .B1(_3159_),
    .Y(_0459_));
 sky130_fd_sc_hd__nand2_1 _4687_ (.A(_3161_),
    .B(_0459_),
    .Y(_0460_));
 sky130_fd_sc_hd__nand3_1 _4688_ (.A(_0456_),
    .B(_0458_),
    .C(_0460_),
    .Y(_0461_));
 sky130_fd_sc_hd__a32oi_2 _4689_ (.A1(_3526_),
    .A2(_3527_),
    .A3(_3525_),
    .B1(_3533_),
    .B2(_0106_),
    .Y(_0462_));
 sky130_fd_sc_hd__o211ai_1 _4690_ (.A1(_3165_),
    .A2(_3164_),
    .B1(_3161_),
    .C1(_3159_),
    .Y(_0463_));
 sky130_fd_sc_hd__nand2_1 _4691_ (.A(_0459_),
    .B(_0457_),
    .Y(_0464_));
 sky130_fd_sc_hd__nand3_2 _4692_ (.A(_0462_),
    .B(_0463_),
    .C(_0464_),
    .Y(_0465_));
 sky130_fd_sc_hd__inv_2 _4693_ (.A(_3516_),
    .Y(_0466_));
 sky130_fd_sc_hd__o21ai_1 _4694_ (.A1(_3346_),
    .A2(_0466_),
    .B1(_3520_),
    .Y(_0467_));
 sky130_fd_sc_hd__nand2_1 _4695_ (.A(_0465_),
    .B(_0467_),
    .Y(_0468_));
 sky130_fd_sc_hd__nand2_1 _4696_ (.A(_0461_),
    .B(_0468_),
    .Y(_0469_));
 sky130_fd_sc_hd__a21o_1 _4697_ (.A1(_3171_),
    .A2(_3168_),
    .B1(_3107_),
    .X(_0470_));
 sky130_fd_sc_hd__nand3_2 _4698_ (.A(_3171_),
    .B(_3168_),
    .C(_3107_),
    .Y(_0471_));
 sky130_fd_sc_hd__nand3_2 _4699_ (.A(_0469_),
    .B(_0470_),
    .C(_0471_),
    .Y(_0472_));
 sky130_fd_sc_hd__a21boi_1 _4700_ (.A1(_0110_),
    .A2(_0112_),
    .B1_N(_0105_),
    .Y(_0473_));
 sky130_fd_sc_hd__a31oi_1 _4701_ (.A1(_3518_),
    .A2(_3519_),
    .A3(_3384_),
    .B1(_3351_),
    .Y(_0474_));
 sky130_fd_sc_hd__o2bb2ai_1 _4702_ (.A1_N(_0465_),
    .A2_N(_0461_),
    .B1(_0474_),
    .B2(_0466_),
    .Y(_0475_));
 sky130_fd_sc_hd__nand3_1 _4703_ (.A(_0465_),
    .B(_0461_),
    .C(_0467_),
    .Y(_0476_));
 sky130_fd_sc_hd__nand3_1 _4704_ (.A(_0473_),
    .B(_0475_),
    .C(_0476_),
    .Y(_0477_));
 sky130_fd_sc_hd__a31o_1 _4705_ (.A1(_0456_),
    .A2(_0458_),
    .A3(_0460_),
    .B1(_0467_),
    .X(_0478_));
 sky130_fd_sc_hd__a22oi_4 _4706_ (.A1(_0465_),
    .A2(_0478_),
    .B1(_0470_),
    .B2(_0471_),
    .Y(_0479_));
 sky130_fd_sc_hd__a21oi_1 _4707_ (.A1(_0472_),
    .A2(_0477_),
    .B1(_0479_),
    .Y(_0480_));
 sky130_fd_sc_hd__a21oi_1 _4708_ (.A1(_0116_),
    .A2(_0454_),
    .B1(_0480_),
    .Y(_0481_));
 sky130_fd_sc_hd__o21ai_4 _4709_ (.A1(_0120_),
    .A2(_0453_),
    .B1(_0481_),
    .Y(_0482_));
 sky130_fd_sc_hd__a21oi_2 _4710_ (.A1(_0475_),
    .A2(_0476_),
    .B1(_0473_),
    .Y(_0483_));
 sky130_fd_sc_hd__o21ai_4 _4711_ (.A1(_0479_),
    .A2(_0483_),
    .B1(_0472_),
    .Y(_0484_));
 sky130_fd_sc_hd__a21o_1 _4712_ (.A1(_3011_),
    .A2(_3175_),
    .B1(_1488_),
    .X(_0485_));
 sky130_fd_sc_hd__o211ai_1 _4713_ (.A1(_3179_),
    .A2(_1477_),
    .B1(_3011_),
    .C1(_3175_),
    .Y(_0486_));
 sky130_fd_sc_hd__nand3_1 _4714_ (.A(_0485_),
    .B(_3172_),
    .C(_0486_),
    .Y(_0487_));
 sky130_fd_sc_hd__and2_2 _4715_ (.A(_3181_),
    .B(_0487_),
    .X(_0488_));
 sky130_fd_sc_hd__nand3_1 _4716_ (.A(_0482_),
    .B(_0484_),
    .C(_0488_),
    .Y(_0489_));
 sky130_fd_sc_hd__o21ai_2 _4717_ (.A1(_3086_),
    .A2(_3084_),
    .B1(_1662_),
    .Y(_0490_));
 sky130_fd_sc_hd__a21o_1 _4718_ (.A1(_3076_),
    .A2(_3082_),
    .B1(_0490_),
    .X(_0491_));
 sky130_fd_sc_hd__nand3_1 _4719_ (.A(_0490_),
    .B(_3076_),
    .C(_3082_),
    .Y(_0492_));
 sky130_fd_sc_hd__nand3_2 _4720_ (.A(_0491_),
    .B(_0492_),
    .C(_3018_),
    .Y(_0493_));
 sky130_fd_sc_hd__nand2_1 _4721_ (.A(_3088_),
    .B(_0493_),
    .Y(_0494_));
 sky130_fd_sc_hd__a21oi_2 _4722_ (.A1(_3181_),
    .A2(_0489_),
    .B1(_0494_),
    .Y(_0495_));
 sky130_fd_sc_hd__nor2_1 _4723_ (.A(_3073_),
    .B(_3074_),
    .Y(_0496_));
 sky130_fd_sc_hd__a21oi_1 _4724_ (.A1(_3062_),
    .A2(_3063_),
    .B1(_3020_),
    .Y(_0497_));
 sky130_fd_sc_hd__a21o_1 _4725_ (.A1(_3064_),
    .A2(_0496_),
    .B1(_0497_),
    .X(_0498_));
 sky130_fd_sc_hd__o2bb2ai_1 _4726_ (.A1_N(net294),
    .A2_N(net103),
    .B1(net309),
    .B2(_1869_),
    .Y(_0499_));
 sky130_fd_sc_hd__nand4_2 _4727_ (.A(_2794_),
    .B(net103),
    .C(net294),
    .D(net98),
    .Y(_0500_));
 sky130_fd_sc_hd__a22oi_2 _4728_ (.A1(net281),
    .A2(net110),
    .B1(_0499_),
    .B2(_0500_),
    .Y(_0501_));
 sky130_fd_sc_hd__and3_1 _4729_ (.A(net98),
    .B(net294),
    .C(net105),
    .X(_0502_));
 sky130_fd_sc_hd__nand2_1 _4730_ (.A(net281),
    .B(net110),
    .Y(_0503_));
 sky130_fd_sc_hd__a22oi_4 _4731_ (.A1(net294),
    .A2(net103),
    .B1(_2794_),
    .B2(net98),
    .Y(_0504_));
 sky130_fd_sc_hd__a211oi_4 _4732_ (.A1(_0502_),
    .A2(_2973_),
    .B1(_0503_),
    .C1(_0504_),
    .Y(_0505_));
 sky130_fd_sc_hd__nand2_1 _4733_ (.A(net295),
    .B(net111),
    .Y(_0506_));
 sky130_fd_sc_hd__o22ai_4 _4734_ (.A1(net320),
    .A2(_3023_),
    .B1(_0506_),
    .B2(_3025_),
    .Y(_0507_));
 sky130_fd_sc_hd__o21bai_4 _4735_ (.A1(_0501_),
    .A2(_0505_),
    .B1_N(_0507_),
    .Y(_0508_));
 sky130_fd_sc_hd__clkbuf_8 _4736_ (.A(_3381_),
    .X(_0509_));
 sky130_fd_sc_hd__o2bb2ai_1 _4737_ (.A1_N(_0499_),
    .A2_N(_0500_),
    .B1(_0509_),
    .B2(_1771_),
    .Y(_0510_));
 sky130_fd_sc_hd__nand4_1 _4738_ (.A(_0499_),
    .B(_0500_),
    .C(net281),
    .D(net110),
    .Y(_0511_));
 sky130_fd_sc_hd__nand3_1 _4739_ (.A(_0510_),
    .B(_0511_),
    .C(_0507_),
    .Y(_0512_));
 sky130_fd_sc_hd__nand4_2 _4740_ (.A(net270),
    .B(net116),
    .C(net253),
    .D(net122),
    .Y(_0513_));
 sky130_fd_sc_hd__a22o_1 _4741_ (.A1(net270),
    .A2(net116),
    .B1(net253),
    .B2(net122),
    .X(_0514_));
 sky130_fd_sc_hd__a22o_1 _4742_ (.A1(net253),
    .A2(net129),
    .B1(_0513_),
    .B2(_0514_),
    .X(_0515_));
 sky130_fd_sc_hd__nand4_2 _4743_ (.A(_0514_),
    .B(net129),
    .C(net253),
    .D(_0513_),
    .Y(_0516_));
 sky130_fd_sc_hd__nand2_2 _4744_ (.A(_0515_),
    .B(_0516_),
    .Y(_0517_));
 sky130_fd_sc_hd__a21o_1 _4745_ (.A1(_0508_),
    .A2(_0512_),
    .B1(_0517_),
    .X(_0518_));
 sky130_fd_sc_hd__nand2_2 _4746_ (.A(_0510_),
    .B(_0507_),
    .Y(_0519_));
 sky130_fd_sc_hd__o211ai_4 _4747_ (.A1(_0505_),
    .A2(_0519_),
    .B1(_0517_),
    .C1(_0508_),
    .Y(_0520_));
 sky130_fd_sc_hd__a21oi_1 _4748_ (.A1(_3026_),
    .A2(_3028_),
    .B1(_3032_),
    .Y(_0521_));
 sky130_fd_sc_hd__o21a_1 _4749_ (.A1(_3038_),
    .A2(_0521_),
    .B1(_3033_),
    .X(_0522_));
 sky130_fd_sc_hd__nand3_2 _4750_ (.A(_0518_),
    .B(_0520_),
    .C(_0522_),
    .Y(_0523_));
 sky130_fd_sc_hd__a21bo_1 _4751_ (.A1(_0508_),
    .A2(_0512_),
    .B1_N(_0517_),
    .X(_0524_));
 sky130_fd_sc_hd__nand4_2 _4752_ (.A(_0508_),
    .B(_0512_),
    .C(_0515_),
    .D(_0516_),
    .Y(_0525_));
 sky130_fd_sc_hd__o21ai_1 _4753_ (.A1(_3038_),
    .A2(_0521_),
    .B1(_3033_),
    .Y(_0526_));
 sky130_fd_sc_hd__nand3_4 _4754_ (.A(_0524_),
    .B(_0525_),
    .C(_0526_),
    .Y(_0527_));
 sky130_fd_sc_hd__nand2_1 _4755_ (.A(_0523_),
    .B(_0527_),
    .Y(_0528_));
 sky130_fd_sc_hd__nor2_1 _4756_ (.A(_2642_),
    .B(_2675_),
    .Y(_0529_));
 sky130_fd_sc_hd__nand2_1 _4757_ (.A(net253),
    .B(net130),
    .Y(_0530_));
 sky130_fd_sc_hd__a22oi_1 _4758_ (.A1(net281),
    .A2(net116),
    .B1(net122),
    .B2(net270),
    .Y(_0531_));
 sky130_fd_sc_hd__o21ai_1 _4759_ (.A1(_0530_),
    .A2(_0531_),
    .B1(_3034_),
    .Y(_0532_));
 sky130_fd_sc_hd__nand2_1 _4760_ (.A(_0529_),
    .B(_0532_),
    .Y(_0533_));
 sky130_fd_sc_hd__a21o_1 _4761_ (.A1(_2577_),
    .A2(_2610_),
    .B1(_0532_),
    .X(_0534_));
 sky130_fd_sc_hd__a21oi_1 _4762_ (.A1(_0533_),
    .A2(_0534_),
    .B1(_3059_),
    .Y(_0535_));
 sky130_fd_sc_hd__and3_1 _4763_ (.A(_0533_),
    .B(_0534_),
    .C(_3059_),
    .X(_0536_));
 sky130_fd_sc_hd__nor2_2 _4764_ (.A(_0535_),
    .B(_0536_),
    .Y(_0537_));
 sky130_fd_sc_hd__nand2_1 _4765_ (.A(_0528_),
    .B(_0537_),
    .Y(_0538_));
 sky130_fd_sc_hd__nand2_1 _4766_ (.A(_3043_),
    .B(_3061_),
    .Y(_0539_));
 sky130_fd_sc_hd__nand2_1 _4767_ (.A(_3048_),
    .B(_0539_),
    .Y(_0540_));
 sky130_fd_sc_hd__o211ai_1 _4768_ (.A1(_0535_),
    .A2(_0536_),
    .B1(_0523_),
    .C1(_0527_),
    .Y(_0541_));
 sky130_fd_sc_hd__nand3_2 _4769_ (.A(_0538_),
    .B(_0540_),
    .C(_0541_),
    .Y(_0542_));
 sky130_fd_sc_hd__a21boi_1 _4770_ (.A1(_3043_),
    .A2(_3061_),
    .B1_N(_3048_),
    .Y(_0543_));
 sky130_fd_sc_hd__nand3_1 _4771_ (.A(_0523_),
    .B(_0527_),
    .C(_0537_),
    .Y(_0544_));
 sky130_fd_sc_hd__o2bb2ai_1 _4772_ (.A1_N(_0523_),
    .A2_N(_0527_),
    .B1(_0535_),
    .B2(_0536_),
    .Y(_0545_));
 sky130_fd_sc_hd__nand3_2 _4773_ (.A(_0543_),
    .B(_0544_),
    .C(_0545_),
    .Y(_0546_));
 sky130_fd_sc_hd__a31o_1 _4774_ (.A1(net260),
    .A2(net144),
    .A3(net137),
    .B1(_2642_),
    .X(_0547_));
 sky130_fd_sc_hd__o311a_1 _4775_ (.A1(_3051_),
    .A2(_3052_),
    .A3(_3053_),
    .B1(_3054_),
    .C1(_0547_),
    .X(_0548_));
 sky130_fd_sc_hd__or3_1 _4776_ (.A(_3086_),
    .B(_3084_),
    .C(_0548_),
    .X(_0549_));
 sky130_fd_sc_hd__o22a_2 _4777_ (.A1(_3086_),
    .A2(_3084_),
    .B1(_3057_),
    .B2(_0548_),
    .X(_0550_));
 sky130_fd_sc_hd__inv_2 _4778_ (.A(_0550_),
    .Y(_0551_));
 sky130_fd_sc_hd__o21ai_1 _4779_ (.A1(_3057_),
    .A2(_0549_),
    .B1(_0551_),
    .Y(_0552_));
 sky130_fd_sc_hd__a21o_1 _4780_ (.A1(_0542_),
    .A2(_0546_),
    .B1(_0552_),
    .X(_0553_));
 sky130_fd_sc_hd__nand3_1 _4781_ (.A(_0552_),
    .B(_0542_),
    .C(_0546_),
    .Y(_0554_));
 sky130_fd_sc_hd__nand3_2 _4782_ (.A(_0498_),
    .B(_0553_),
    .C(_0554_),
    .Y(_0555_));
 sky130_fd_sc_hd__a21oi_1 _4783_ (.A1(_3064_),
    .A2(_0496_),
    .B1(_0497_),
    .Y(_0556_));
 sky130_fd_sc_hd__o21a_1 _4784_ (.A1(_3057_),
    .A2(_0549_),
    .B1(_0551_),
    .X(_0557_));
 sky130_fd_sc_hd__a21o_1 _4785_ (.A1(_0542_),
    .A2(_0546_),
    .B1(_0557_),
    .X(_0558_));
 sky130_fd_sc_hd__o2111ai_2 _4786_ (.A1(_0549_),
    .A2(_3057_),
    .B1(_0551_),
    .C1(_0542_),
    .D1(_0546_),
    .Y(_0559_));
 sky130_fd_sc_hd__nand3_1 _4787_ (.A(_0556_),
    .B(_0558_),
    .C(_0559_),
    .Y(_0560_));
 sky130_fd_sc_hd__a2bb2o_1 _4788_ (.A1_N(_3179_),
    .A2_N(_3069_),
    .B1(_0555_),
    .B2(_0560_),
    .X(_0561_));
 sky130_fd_sc_hd__and3_1 _4789_ (.A(_0542_),
    .B(_0546_),
    .C(_0557_),
    .X(_0562_));
 sky130_fd_sc_hd__nand2_1 _4790_ (.A(_0556_),
    .B(_0558_),
    .Y(_0563_));
 sky130_fd_sc_hd__o211ai_1 _4791_ (.A1(_0562_),
    .A2(_0563_),
    .B1(_0555_),
    .C1(_3071_),
    .Y(_0564_));
 sky130_fd_sc_hd__o211a_1 _4792_ (.A1(_2945_),
    .A2(_3079_),
    .B1(_3080_),
    .C1(_3081_),
    .X(_0565_));
 sky130_fd_sc_hd__a21oi_1 _4793_ (.A1(_0490_),
    .A2(_3076_),
    .B1(_0565_),
    .Y(_0566_));
 sky130_fd_sc_hd__nand3_2 _4794_ (.A(_0561_),
    .B(_0564_),
    .C(_0566_),
    .Y(_0567_));
 sky130_fd_sc_hd__a21o_1 _4795_ (.A1(_0490_),
    .A2(_3076_),
    .B1(_0565_),
    .X(_0568_));
 sky130_fd_sc_hd__o221ai_1 _4796_ (.A1(_3179_),
    .A2(_3069_),
    .B1(_0562_),
    .B2(_0563_),
    .C1(_0555_),
    .Y(_0569_));
 sky130_fd_sc_hd__nand2_1 _4797_ (.A(_0555_),
    .B(_0560_),
    .Y(_0570_));
 sky130_fd_sc_hd__nand2_1 _4798_ (.A(_0570_),
    .B(_3071_),
    .Y(_0571_));
 sky130_fd_sc_hd__nand3_1 _4799_ (.A(_0568_),
    .B(_0569_),
    .C(_0571_),
    .Y(_0572_));
 sky130_fd_sc_hd__nand2_1 _4800_ (.A(_0567_),
    .B(_0572_),
    .Y(_0573_));
 sky130_fd_sc_hd__o21bai_1 _4801_ (.A1(_3089_),
    .A2(_0495_),
    .B1_N(_0573_),
    .Y(_0574_));
 sky130_fd_sc_hd__a211o_1 _4802_ (.A1(_0567_),
    .A2(_0572_),
    .B1(_3089_),
    .C1(_0495_),
    .X(_0575_));
 sky130_fd_sc_hd__and2_1 _4803_ (.A(_0574_),
    .B(_0575_),
    .X(_0576_));
 sky130_fd_sc_hd__clkbuf_1 _4804_ (.A(_0576_),
    .X(_0076_));
 sky130_fd_sc_hd__a21bo_1 _4805_ (.A1(_0557_),
    .A2(_0546_),
    .B1_N(_0542_),
    .X(_0577_));
 sky130_fd_sc_hd__o21a_1 _4806_ (.A1(net116),
    .A2(net122),
    .B1(net252),
    .X(_0578_));
 sky130_fd_sc_hd__nand3_2 _4807_ (.A(net116),
    .B(net252),
    .C(net122),
    .Y(_0579_));
 sky130_fd_sc_hd__and4_2 _4808_ (.A(_0578_),
    .B(net129),
    .C(net252),
    .D(_0579_),
    .X(_0580_));
 sky130_fd_sc_hd__o2bb2a_2 _4809_ (.A1_N(_0579_),
    .A2_N(_0578_),
    .B1(_1423_),
    .B2(_2931_),
    .X(_0581_));
 sky130_fd_sc_hd__nand3_1 _4810_ (.A(net97),
    .B(net103),
    .C(net281),
    .Y(_0582_));
 sky130_fd_sc_hd__nor2_1 _4811_ (.A(net294),
    .B(_0582_),
    .Y(_0583_));
 sky130_fd_sc_hd__a22oi_2 _4812_ (.A1(net104),
    .A2(net281),
    .B1(_3021_),
    .B2(net98),
    .Y(_0584_));
 sky130_fd_sc_hd__o22ai_2 _4813_ (.A1(_1771_),
    .A2(_2928_),
    .B1(_0583_),
    .B2(_0584_),
    .Y(_0585_));
 sky130_fd_sc_hd__o2bb2ai_1 _4814_ (.A1_N(net105),
    .A2_N(net281),
    .B1(net294),
    .B2(_1869_),
    .Y(_0586_));
 sky130_fd_sc_hd__o2111ai_2 _4815_ (.A1(net294),
    .A2(_0582_),
    .B1(net269),
    .C1(net110),
    .D1(_0586_),
    .Y(_0587_));
 sky130_fd_sc_hd__o21ai_2 _4816_ (.A1(_0503_),
    .A2(_0504_),
    .B1(_0500_),
    .Y(_0588_));
 sky130_fd_sc_hd__a21oi_1 _4817_ (.A1(_0585_),
    .A2(_0587_),
    .B1(_0588_),
    .Y(_0589_));
 sky130_fd_sc_hd__nand4_1 _4818_ (.A(_3022_),
    .B(net104),
    .C(net281),
    .D(net98),
    .Y(_0590_));
 sky130_fd_sc_hd__nand3_1 _4819_ (.A(_0586_),
    .B(net269),
    .C(_0590_),
    .Y(_0591_));
 sky130_fd_sc_hd__o211a_2 _4820_ (.A1(_2920_),
    .A2(_0591_),
    .B1(_0588_),
    .C1(_0585_),
    .X(_0592_));
 sky130_fd_sc_hd__o22ai_4 _4821_ (.A1(_0580_),
    .A2(_0581_),
    .B1(_0589_),
    .B2(_0592_),
    .Y(_0593_));
 sky130_fd_sc_hd__a21o_1 _4822_ (.A1(_0585_),
    .A2(_0587_),
    .B1(_0588_),
    .X(_0594_));
 sky130_fd_sc_hd__o211ai_1 _4823_ (.A1(_2920_),
    .A2(_0591_),
    .B1(_0588_),
    .C1(_0585_),
    .Y(_0595_));
 sky130_fd_sc_hd__nor2_2 _4824_ (.A(_0580_),
    .B(_0581_),
    .Y(_0596_));
 sky130_fd_sc_hd__nand3_1 _4825_ (.A(_0594_),
    .B(_0595_),
    .C(_0596_),
    .Y(_0597_));
 sky130_fd_sc_hd__a21oi_1 _4826_ (.A1(_0510_),
    .A2(_0511_),
    .B1(_0507_),
    .Y(_0598_));
 sky130_fd_sc_hd__o22ai_4 _4827_ (.A1(_0505_),
    .A2(_0519_),
    .B1(_0517_),
    .B2(_0598_),
    .Y(_0599_));
 sky130_fd_sc_hd__a21oi_2 _4828_ (.A1(_0593_),
    .A2(_0597_),
    .B1(_0599_),
    .Y(_0600_));
 sky130_fd_sc_hd__nand2_1 _4829_ (.A(_0594_),
    .B(_0596_),
    .Y(_0601_));
 sky130_fd_sc_hd__o211a_1 _4830_ (.A1(_0592_),
    .A2(_0601_),
    .B1(_0599_),
    .C1(_0593_),
    .X(_0602_));
 sky130_fd_sc_hd__o21ai_1 _4831_ (.A1(_3342_),
    .A2(_2931_),
    .B1(_0513_),
    .Y(_0603_));
 sky130_fd_sc_hd__nand2_1 _4832_ (.A(_0514_),
    .B(_0603_),
    .Y(_0604_));
 sky130_fd_sc_hd__o21ai_1 _4833_ (.A1(_2653_),
    .A2(_2675_),
    .B1(_0604_),
    .Y(_0605_));
 sky130_fd_sc_hd__nand4_1 _4834_ (.A(_2577_),
    .B(_2610_),
    .C(_0514_),
    .D(_0603_),
    .Y(_0606_));
 sky130_fd_sc_hd__nand2_1 _4835_ (.A(_0605_),
    .B(_0606_),
    .Y(_0607_));
 sky130_fd_sc_hd__xor2_2 _4836_ (.A(_3059_),
    .B(_0607_),
    .X(_0608_));
 sky130_fd_sc_hd__o21bai_2 _4837_ (.A1(_0600_),
    .A2(_0602_),
    .B1_N(_0608_),
    .Y(_0609_));
 sky130_fd_sc_hd__a21o_1 _4838_ (.A1(_0593_),
    .A2(_0597_),
    .B1(_0599_),
    .X(_0610_));
 sky130_fd_sc_hd__o211ai_1 _4839_ (.A1(_0592_),
    .A2(_0601_),
    .B1(_0599_),
    .C1(_0593_),
    .Y(_0611_));
 sky130_fd_sc_hd__nand3_1 _4840_ (.A(_0610_),
    .B(_0611_),
    .C(_0608_),
    .Y(_0612_));
 sky130_fd_sc_hd__a32oi_4 _4841_ (.A1(_0518_),
    .A2(_0520_),
    .A3(_0522_),
    .B1(_0527_),
    .B2(_0537_),
    .Y(_0613_));
 sky130_fd_sc_hd__a21oi_2 _4842_ (.A1(_0609_),
    .A2(_0612_),
    .B1(_0613_),
    .Y(_0614_));
 sky130_fd_sc_hd__nand2_1 _4843_ (.A(_0608_),
    .B(_0611_),
    .Y(_0615_));
 sky130_fd_sc_hd__o211a_1 _4844_ (.A1(_0600_),
    .A2(_0615_),
    .B1(_0609_),
    .C1(_0613_),
    .X(_0616_));
 sky130_fd_sc_hd__a21boi_1 _4845_ (.A1(_0547_),
    .A2(_0534_),
    .B1_N(_0533_),
    .Y(_0617_));
 sky130_fd_sc_hd__a21oi_1 _4846_ (.A1(_1156_),
    .A2(_1183_),
    .B1(_0617_),
    .Y(_0618_));
 sky130_fd_sc_hd__and3_1 _4847_ (.A(_0617_),
    .B(_1156_),
    .C(_1183_),
    .X(_0619_));
 sky130_fd_sc_hd__or2_1 _4848_ (.A(_0618_),
    .B(_0619_),
    .X(_0620_));
 sky130_fd_sc_hd__clkbuf_2 _4849_ (.A(_0620_),
    .X(_0621_));
 sky130_fd_sc_hd__o21ai_1 _4850_ (.A1(_0614_),
    .A2(_0616_),
    .B1(_0621_),
    .Y(_0622_));
 sky130_fd_sc_hd__o211ai_4 _4851_ (.A1(_0600_),
    .A2(_0615_),
    .B1(_0609_),
    .C1(_0613_),
    .Y(_0623_));
 sky130_fd_sc_hd__inv_2 _4852_ (.A(_0621_),
    .Y(_0624_));
 sky130_fd_sc_hd__nand3b_1 _4853_ (.A_N(_0614_),
    .B(_0623_),
    .C(_0624_),
    .Y(_0625_));
 sky130_fd_sc_hd__nand3_2 _4854_ (.A(_0577_),
    .B(_0622_),
    .C(_0625_),
    .Y(_0626_));
 sky130_fd_sc_hd__a32o_1 _4855_ (.A1(_0543_),
    .A2(_0544_),
    .A3(_0545_),
    .B1(_0542_),
    .B2(_0552_),
    .X(_0627_));
 sky130_fd_sc_hd__nand3b_1 _4856_ (.A_N(_0614_),
    .B(_0623_),
    .C(_0621_),
    .Y(_0628_));
 sky130_fd_sc_hd__o21bai_1 _4857_ (.A1(_0614_),
    .A2(_0616_),
    .B1_N(_0621_),
    .Y(_0629_));
 sky130_fd_sc_hd__nand3_2 _4858_ (.A(_0627_),
    .B(_0628_),
    .C(_0629_),
    .Y(_0630_));
 sky130_fd_sc_hd__nand2_2 _4859_ (.A(_0626_),
    .B(_0630_),
    .Y(_0631_));
 sky130_fd_sc_hd__o2bb2ai_1 _4860_ (.A1_N(_3071_),
    .A2_N(_0555_),
    .B1(_0563_),
    .B2(_0562_),
    .Y(_0632_));
 sky130_fd_sc_hd__a21oi_1 _4861_ (.A1(_0631_),
    .A2(_0550_),
    .B1(_0632_),
    .Y(_0633_));
 sky130_fd_sc_hd__o21ai_2 _4862_ (.A1(_0550_),
    .A2(_0631_),
    .B1(_0633_),
    .Y(_0634_));
 sky130_fd_sc_hd__inv_2 _4863_ (.A(_0634_),
    .Y(_0635_));
 sky130_fd_sc_hd__nand3_1 _4864_ (.A(_0626_),
    .B(_0630_),
    .C(_0550_),
    .Y(_0636_));
 sky130_fd_sc_hd__nand2_1 _4865_ (.A(_0632_),
    .B(_0636_),
    .Y(_0637_));
 sky130_fd_sc_hd__a21o_1 _4866_ (.A1(_0551_),
    .A2(_0631_),
    .B1(_0637_),
    .X(_0638_));
 sky130_fd_sc_hd__inv_2 _4867_ (.A(_0638_),
    .Y(_0639_));
 sky130_fd_sc_hd__o2bb2ai_1 _4868_ (.A1_N(_0567_),
    .A2_N(_0574_),
    .B1(_0635_),
    .B2(_0639_),
    .Y(_0640_));
 sky130_fd_sc_hd__a21oi_1 _4869_ (.A1(_0626_),
    .A2(_0630_),
    .B1(_0550_),
    .Y(_0641_));
 sky130_fd_sc_hd__o2111ai_1 _4870_ (.A1(_0641_),
    .A2(_0637_),
    .B1(_0634_),
    .C1(_0567_),
    .D1(_0574_),
    .Y(_0642_));
 sky130_fd_sc_hd__nand2_1 _4871_ (.A(_0640_),
    .B(_0642_),
    .Y(_0077_));
 sky130_fd_sc_hd__and3_1 _4872_ (.A(_0551_),
    .B(_0626_),
    .C(_0630_),
    .X(_0643_));
 sky130_fd_sc_hd__a31oi_1 _4873_ (.A1(_0556_),
    .A2(_0558_),
    .A3(_0559_),
    .B1(_3071_),
    .Y(_0644_));
 sky130_fd_sc_hd__and3_1 _4874_ (.A(_0498_),
    .B(_0553_),
    .C(_0554_),
    .X(_0645_));
 sky130_fd_sc_hd__o2bb2ai_1 _4875_ (.A1_N(_0550_),
    .A2_N(_0631_),
    .B1(_0644_),
    .B2(_0645_),
    .Y(_0646_));
 sky130_fd_sc_hd__o22ai_2 _4876_ (.A1(_0641_),
    .A2(_0637_),
    .B1(_0643_),
    .B2(_0646_),
    .Y(_0647_));
 sky130_fd_sc_hd__nand4_1 _4877_ (.A(_3088_),
    .B(_3181_),
    .C(_0487_),
    .D(_0493_),
    .Y(_0648_));
 sky130_fd_sc_hd__nor3_1 _4878_ (.A(_0573_),
    .B(_0647_),
    .C(_0648_),
    .Y(_0649_));
 sky130_fd_sc_hd__nand3_1 _4879_ (.A(_0482_),
    .B(_0649_),
    .C(_0484_),
    .Y(_0650_));
 sky130_fd_sc_hd__nor2_1 _4880_ (.A(_0573_),
    .B(_0647_),
    .Y(_0651_));
 sky130_fd_sc_hd__a32oi_1 _4881_ (.A1(_3018_),
    .A2(_0491_),
    .A3(_0492_),
    .B1(_3088_),
    .B2(_3181_),
    .Y(_0652_));
 sky130_fd_sc_hd__a21boi_1 _4882_ (.A1(_0567_),
    .A2(_0638_),
    .B1_N(_0634_),
    .Y(_0653_));
 sky130_fd_sc_hd__a21oi_1 _4883_ (.A1(_0651_),
    .A2(_0652_),
    .B1(_0653_),
    .Y(_0654_));
 sky130_fd_sc_hd__nand2_1 _4884_ (.A(_0650_),
    .B(_0654_),
    .Y(_0655_));
 sky130_fd_sc_hd__nand4_2 _4885_ (.A(_0578_),
    .B(net129),
    .C(net252),
    .D(_0579_),
    .Y(_0656_));
 sky130_fd_sc_hd__a211o_1 _4886_ (.A1(_0579_),
    .A2(_0656_),
    .B1(_2653_),
    .C1(_2675_),
    .X(_0657_));
 sky130_fd_sc_hd__and3_1 _4887_ (.A(net116),
    .B(net252),
    .C(net122),
    .X(_0658_));
 sky130_fd_sc_hd__a31o_1 _4888_ (.A1(_0578_),
    .A2(net129),
    .A3(net252),
    .B1(_0658_),
    .X(_0659_));
 sky130_fd_sc_hd__o22a_1 _4889_ (.A1(_2599_),
    .A2(_2653_),
    .B1(_0659_),
    .B2(_0529_),
    .X(_0660_));
 sky130_fd_sc_hd__a21o_1 _4890_ (.A1(_2577_),
    .A2(_2610_),
    .B1(_0659_),
    .X(_0661_));
 sky130_fd_sc_hd__a21oi_1 _4891_ (.A1(_0657_),
    .A2(_0661_),
    .B1(_0547_),
    .Y(_0662_));
 sky130_fd_sc_hd__a21oi_2 _4892_ (.A1(_0657_),
    .A2(_0660_),
    .B1(_0662_),
    .Y(_0663_));
 sky130_fd_sc_hd__clkbuf_2 _4893_ (.A(_0663_),
    .X(_0664_));
 sky130_fd_sc_hd__o2bb2ai_1 _4894_ (.A1_N(net103),
    .A2_N(net269),
    .B1(net286),
    .B2(_3127_),
    .Y(_0665_));
 sky130_fd_sc_hd__nand4_2 _4895_ (.A(_3381_),
    .B(net269),
    .C(net97),
    .D(net103),
    .Y(_0666_));
 sky130_fd_sc_hd__nand2_1 _4896_ (.A(net110),
    .B(net252),
    .Y(_0667_));
 sky130_fd_sc_hd__a21o_1 _4897_ (.A1(_0665_),
    .A2(_0666_),
    .B1(_0667_),
    .X(_0668_));
 sky130_fd_sc_hd__o211ai_1 _4898_ (.A1(_2920_),
    .A2(_3176_),
    .B1(_0665_),
    .C1(_0666_),
    .Y(_0669_));
 sky130_fd_sc_hd__nor2_1 _4899_ (.A(_2920_),
    .B(_2929_),
    .Y(_0670_));
 sky130_fd_sc_hd__a21oi_1 _4900_ (.A1(_0586_),
    .A2(_0670_),
    .B1(_0583_),
    .Y(_0671_));
 sky130_fd_sc_hd__nand3_1 _4901_ (.A(_0668_),
    .B(_0669_),
    .C(_0671_),
    .Y(_0672_));
 sky130_fd_sc_hd__a41o_1 _4902_ (.A1(_0509_),
    .A2(net269),
    .A3(net97),
    .A4(net103),
    .B1(_0667_),
    .X(_0673_));
 sky130_fd_sc_hd__a22oi_4 _4903_ (.A1(net103),
    .A2(net269),
    .B1(_0509_),
    .B2(net97),
    .Y(_0674_));
 sky130_fd_sc_hd__nand2_1 _4904_ (.A(net110),
    .B(net269),
    .Y(_0675_));
 sky130_fd_sc_hd__o21ai_1 _4905_ (.A1(_0675_),
    .A2(_0584_),
    .B1(_0590_),
    .Y(_0676_));
 sky130_fd_sc_hd__o2bb2ai_1 _4906_ (.A1_N(_0665_),
    .A2_N(_0666_),
    .B1(_2920_),
    .B2(_3176_),
    .Y(_0677_));
 sky130_fd_sc_hd__o211ai_4 _4907_ (.A1(_0673_),
    .A2(_0674_),
    .B1(_0676_),
    .C1(_0677_),
    .Y(_0678_));
 sky130_fd_sc_hd__nand2_1 _4908_ (.A(_0672_),
    .B(_0678_),
    .Y(_0679_));
 sky130_fd_sc_hd__nand2_1 _4909_ (.A(_0679_),
    .B(_0596_),
    .Y(_0680_));
 sky130_fd_sc_hd__a21oi_1 _4910_ (.A1(_0594_),
    .A2(_0596_),
    .B1(_0592_),
    .Y(_0681_));
 sky130_fd_sc_hd__o211ai_2 _4911_ (.A1(_0580_),
    .A2(_0581_),
    .B1(_0672_),
    .C1(_0678_),
    .Y(_0682_));
 sky130_fd_sc_hd__nand3_1 _4912_ (.A(_0680_),
    .B(_0681_),
    .C(_0682_),
    .Y(_0683_));
 sky130_fd_sc_hd__a21oi_1 _4913_ (.A1(_0682_),
    .A2(_0680_),
    .B1(_0681_),
    .Y(_0684_));
 sky130_fd_sc_hd__a21oi_1 _4914_ (.A1(_0663_),
    .A2(_0683_),
    .B1(_0684_),
    .Y(_0685_));
 sky130_fd_sc_hd__o21ai_1 _4915_ (.A1(_0664_),
    .A2(_0683_),
    .B1(_0685_),
    .Y(_0686_));
 sky130_fd_sc_hd__a21oi_1 _4916_ (.A1(_0610_),
    .A2(_0608_),
    .B1(_0602_),
    .Y(_0687_));
 sky130_fd_sc_hd__nand2_1 _4917_ (.A(_0664_),
    .B(_0684_),
    .Y(_0688_));
 sky130_fd_sc_hd__nand3_1 _4918_ (.A(_0686_),
    .B(_0687_),
    .C(_0688_),
    .Y(_0689_));
 sky130_fd_sc_hd__a21o_1 _4919_ (.A1(_0610_),
    .A2(_0608_),
    .B1(_0602_),
    .X(_0690_));
 sky130_fd_sc_hd__and3_1 _4920_ (.A(_0680_),
    .B(_0681_),
    .C(_0682_),
    .X(_0691_));
 sky130_fd_sc_hd__o21bai_1 _4921_ (.A1(_0684_),
    .A2(_0691_),
    .B1_N(_0663_),
    .Y(_0692_));
 sky130_fd_sc_hd__nand3b_1 _4922_ (.A_N(_0684_),
    .B(_0683_),
    .C(_0664_),
    .Y(_0693_));
 sky130_fd_sc_hd__nand3_1 _4923_ (.A(_0690_),
    .B(_0692_),
    .C(_0693_),
    .Y(_0694_));
 sky130_fd_sc_hd__o32a_1 _4924_ (.A1(_2653_),
    .A2(_2675_),
    .A3(_0604_),
    .B1(_3059_),
    .B2(_0607_),
    .X(_0695_));
 sky130_fd_sc_hd__a21oi_1 _4925_ (.A1(_1165_),
    .A2(_1193_),
    .B1(_0695_),
    .Y(_0696_));
 sky130_fd_sc_hd__and3_1 _4926_ (.A(_0695_),
    .B(_1165_),
    .C(_1193_),
    .X(_0697_));
 sky130_fd_sc_hd__or2_1 _4927_ (.A(_0696_),
    .B(_0697_),
    .X(_0698_));
 sky130_fd_sc_hd__nand3_1 _4928_ (.A(_0689_),
    .B(_0694_),
    .C(_0698_),
    .Y(_0699_));
 sky130_fd_sc_hd__a21o_1 _4929_ (.A1(_0689_),
    .A2(_0694_),
    .B1(_0698_),
    .X(_0700_));
 sky130_fd_sc_hd__nand2_1 _4930_ (.A(_0699_),
    .B(_0700_),
    .Y(_0701_));
 sky130_fd_sc_hd__o21ai_1 _4931_ (.A1(_0621_),
    .A2(_0614_),
    .B1(_0623_),
    .Y(_0702_));
 sky130_fd_sc_hd__nand2_1 _4932_ (.A(_0701_),
    .B(_0702_),
    .Y(_0703_));
 sky130_fd_sc_hd__o211ai_1 _4933_ (.A1(_0616_),
    .A2(_0701_),
    .B1(_0618_),
    .C1(_0703_),
    .Y(_0704_));
 sky130_fd_sc_hd__o2111ai_2 _4934_ (.A1(_0621_),
    .A2(_0614_),
    .B1(_0623_),
    .C1(_0699_),
    .D1(_0700_),
    .Y(_0705_));
 sky130_fd_sc_hd__a21o_1 _4935_ (.A1(_0703_),
    .A2(_0705_),
    .B1(_0618_),
    .X(_0706_));
 sky130_fd_sc_hd__o21ai_1 _4936_ (.A1(_0551_),
    .A2(_0631_),
    .B1(_0626_),
    .Y(_0707_));
 sky130_fd_sc_hd__a21oi_1 _4937_ (.A1(_0704_),
    .A2(_0706_),
    .B1(_0707_),
    .Y(_0708_));
 sky130_fd_sc_hd__nand3_1 _4938_ (.A(_0707_),
    .B(_0704_),
    .C(_0706_),
    .Y(_0709_));
 sky130_fd_sc_hd__or2b_1 _4939_ (.A(_0708_),
    .B_N(_0709_),
    .X(_0710_));
 sky130_fd_sc_hd__xnor2_1 _4940_ (.A(_0655_),
    .B(_0710_),
    .Y(_0078_));
 sky130_fd_sc_hd__a21boi_1 _4941_ (.A1(_0618_),
    .A2(_0705_),
    .B1_N(_0703_),
    .Y(_0711_));
 sky130_fd_sc_hd__o21a_1 _4942_ (.A1(net104),
    .A2(net110),
    .B1(net255),
    .X(_0712_));
 sky130_fd_sc_hd__nand3_2 _4943_ (.A(net104),
    .B(net110),
    .C(net255),
    .Y(_0713_));
 sky130_fd_sc_hd__a22o_1 _4944_ (.A1(net97),
    .A2(_2929_),
    .B1(_0712_),
    .B2(_0713_),
    .X(_0714_));
 sky130_fd_sc_hd__nand4_1 _4945_ (.A(_2929_),
    .B(_0712_),
    .C(_0713_),
    .D(net97),
    .Y(_0715_));
 sky130_fd_sc_hd__o21ai_2 _4946_ (.A1(_0667_),
    .A2(_0674_),
    .B1(_0666_),
    .Y(_0716_));
 sky130_fd_sc_hd__a21oi_2 _4947_ (.A1(_0714_),
    .A2(_0715_),
    .B1(_0716_),
    .Y(_0717_));
 sky130_fd_sc_hd__o211a_1 _4948_ (.A1(_3127_),
    .A2(net269),
    .B1(_0713_),
    .C1(_0712_),
    .X(_0718_));
 sky130_fd_sc_hd__nand2_1 _4949_ (.A(_2929_),
    .B(net97),
    .Y(_0719_));
 sky130_fd_sc_hd__a21oi_1 _4950_ (.A1(_0712_),
    .A2(_0713_),
    .B1(_0719_),
    .Y(_0720_));
 sky130_fd_sc_hd__o21a_1 _4951_ (.A1(_0718_),
    .A2(_0720_),
    .B1(_0716_),
    .X(_0721_));
 sky130_fd_sc_hd__a22o_1 _4952_ (.A1(net252),
    .A2(net129),
    .B1(_0579_),
    .B2(_0578_),
    .X(_0722_));
 sky130_fd_sc_hd__nand2_2 _4953_ (.A(_0656_),
    .B(_0722_),
    .Y(_0723_));
 sky130_fd_sc_hd__o21ai_1 _4954_ (.A1(_0717_),
    .A2(_0721_),
    .B1(_0723_),
    .Y(_0724_));
 sky130_fd_sc_hd__a21o_1 _4955_ (.A1(_0714_),
    .A2(_0715_),
    .B1(_0716_),
    .X(_0725_));
 sky130_fd_sc_hd__o21ai_2 _4956_ (.A1(_0718_),
    .A2(_0720_),
    .B1(_0716_),
    .Y(_0726_));
 sky130_fd_sc_hd__nand3_1 _4957_ (.A(_0725_),
    .B(_0726_),
    .C(_0596_),
    .Y(_0727_));
 sky130_fd_sc_hd__o211a_1 _4958_ (.A1(_0582_),
    .A2(net294),
    .B1(_0669_),
    .C1(_0587_),
    .X(_0728_));
 sky130_fd_sc_hd__a22oi_2 _4959_ (.A1(_0728_),
    .A2(_0668_),
    .B1(_0723_),
    .B2(_0678_),
    .Y(_0729_));
 sky130_fd_sc_hd__a21o_1 _4960_ (.A1(_0724_),
    .A2(_0727_),
    .B1(_0729_),
    .X(_0730_));
 sky130_fd_sc_hd__nand3_2 _4961_ (.A(_0729_),
    .B(_0727_),
    .C(_0724_),
    .Y(_0731_));
 sky130_fd_sc_hd__a21o_1 _4962_ (.A1(_0730_),
    .A2(_0731_),
    .B1(_0663_),
    .X(_0732_));
 sky130_fd_sc_hd__nand3_2 _4963_ (.A(_0730_),
    .B(_0731_),
    .C(_0664_),
    .Y(_0733_));
 sky130_fd_sc_hd__a21bo_1 _4964_ (.A1(_0732_),
    .A2(_0733_),
    .B1_N(_0685_),
    .X(_0734_));
 sky130_fd_sc_hd__nand3b_1 _4965_ (.A_N(_0685_),
    .B(_0732_),
    .C(_0733_),
    .Y(_0735_));
 sky130_fd_sc_hd__a2bb2o_1 _4966_ (.A1_N(_0659_),
    .A2_N(_0529_),
    .B1(_2577_),
    .B2(_2664_),
    .X(_0736_));
 sky130_fd_sc_hd__o2bb2a_2 _4967_ (.A1_N(_0657_),
    .A2_N(_0736_),
    .B1(_3086_),
    .B2(_3084_),
    .X(_0737_));
 sky130_fd_sc_hd__and3_1 _4968_ (.A(_0736_),
    .B(_3179_),
    .C(_0657_),
    .X(_0738_));
 sky130_fd_sc_hd__or2_1 _4969_ (.A(_0737_),
    .B(_0738_),
    .X(_0739_));
 sky130_fd_sc_hd__a21o_1 _4970_ (.A1(_0734_),
    .A2(_0735_),
    .B1(_0739_),
    .X(_0740_));
 sky130_fd_sc_hd__a21bo_1 _4971_ (.A1(_0694_),
    .A2(_0698_),
    .B1_N(_0689_),
    .X(_0741_));
 sky130_fd_sc_hd__o211ai_1 _4972_ (.A1(_0737_),
    .A2(_0738_),
    .B1(_0734_),
    .C1(_0735_),
    .Y(_0742_));
 sky130_fd_sc_hd__nand3_1 _4973_ (.A(_0740_),
    .B(_0741_),
    .C(_0742_),
    .Y(_0743_));
 sky130_fd_sc_hd__a21o_1 _4974_ (.A1(_0742_),
    .A2(_0740_),
    .B1(_0741_),
    .X(_0744_));
 sky130_fd_sc_hd__o211ai_1 _4975_ (.A1(_3179_),
    .A2(_0695_),
    .B1(_0743_),
    .C1(_0744_),
    .Y(_0745_));
 sky130_fd_sc_hd__a21bo_1 _4976_ (.A1(_0743_),
    .A2(_0744_),
    .B1_N(_0696_),
    .X(_0746_));
 sky130_fd_sc_hd__nand3_1 _4977_ (.A(_0711_),
    .B(_0745_),
    .C(_0746_),
    .Y(_0747_));
 sky130_fd_sc_hd__a21o_1 _4978_ (.A1(_0745_),
    .A2(_0746_),
    .B1(_0711_),
    .X(_0748_));
 sky130_fd_sc_hd__nand2_1 _4979_ (.A(_0747_),
    .B(_0748_),
    .Y(_0749_));
 sky130_fd_sc_hd__a31o_1 _4980_ (.A1(_0650_),
    .A2(_0654_),
    .A3(_0709_),
    .B1(_0708_),
    .X(_0750_));
 sky130_fd_sc_hd__xor2_1 _4981_ (.A(_0749_),
    .B(_0750_),
    .X(_0079_));
 sky130_fd_sc_hd__a31o_1 _4982_ (.A1(_0656_),
    .A2(_0722_),
    .A3(_0725_),
    .B1(_0721_),
    .X(_0751_));
 sky130_fd_sc_hd__nand3_1 _4983_ (.A(_0713_),
    .B(net97),
    .C(_2929_),
    .Y(_0752_));
 sky130_fd_sc_hd__o2bb2a_1 _4984_ (.A1_N(_0752_),
    .A2_N(_0712_),
    .B1(net255),
    .B2(_3127_),
    .X(_0753_));
 sky130_fd_sc_hd__o21a_2 _4985_ (.A1(_0580_),
    .A2(_0581_),
    .B1(_0753_),
    .X(_0754_));
 sky130_fd_sc_hd__nor2_1 _4986_ (.A(_0753_),
    .B(_0723_),
    .Y(_0755_));
 sky130_fd_sc_hd__nor2_1 _4987_ (.A(_0754_),
    .B(_0755_),
    .Y(_0756_));
 sky130_fd_sc_hd__nand2_1 _4988_ (.A(_0751_),
    .B(_0756_),
    .Y(_0757_));
 sky130_fd_sc_hd__o221ai_4 _4989_ (.A1(_0723_),
    .A2(_0717_),
    .B1(_0754_),
    .B2(_0755_),
    .C1(_0726_),
    .Y(_0758_));
 sky130_fd_sc_hd__and3_1 _4990_ (.A(_0757_),
    .B(_0664_),
    .C(_0758_),
    .X(_0759_));
 sky130_fd_sc_hd__a21oi_1 _4991_ (.A1(_0758_),
    .A2(_0757_),
    .B1(_0664_),
    .Y(_0760_));
 sky130_fd_sc_hd__a211o_1 _4992_ (.A1(_0731_),
    .A2(_0733_),
    .B1(_0759_),
    .C1(_0760_),
    .X(_0761_));
 sky130_fd_sc_hd__o211ai_2 _4993_ (.A1(_0759_),
    .A2(_0760_),
    .B1(_0731_),
    .C1(_0733_),
    .Y(_0762_));
 sky130_fd_sc_hd__a211o_1 _4994_ (.A1(_0761_),
    .A2(_0762_),
    .B1(_0737_),
    .C1(_0738_),
    .X(_0763_));
 sky130_fd_sc_hd__buf_6 _4995_ (.A(_0737_),
    .X(_0764_));
 sky130_fd_sc_hd__o211ai_1 _4996_ (.A1(_0764_),
    .A2(_0738_),
    .B1(_0761_),
    .C1(_0762_),
    .Y(_0765_));
 sky130_fd_sc_hd__nor2_1 _4997_ (.A(_0737_),
    .B(_0738_),
    .Y(_0766_));
 sky130_fd_sc_hd__a21bo_1 _4998_ (.A1(_0734_),
    .A2(_0766_),
    .B1_N(_0735_),
    .X(_0767_));
 sky130_fd_sc_hd__a21boi_1 _4999_ (.A1(_0763_),
    .A2(_0765_),
    .B1_N(_0767_),
    .Y(_0768_));
 sky130_fd_sc_hd__nand3b_1 _5000_ (.A_N(_0767_),
    .B(_0763_),
    .C(_0765_),
    .Y(_0769_));
 sky130_fd_sc_hd__and3b_1 _5001_ (.A_N(_0768_),
    .B(_0769_),
    .C(_0764_),
    .X(_0770_));
 sky130_fd_sc_hd__and2b_1 _5002_ (.A_N(_0768_),
    .B(_0769_),
    .X(_0771_));
 sky130_fd_sc_hd__a21boi_1 _5003_ (.A1(_0696_),
    .A2(_0743_),
    .B1_N(_0744_),
    .Y(_0772_));
 sky130_fd_sc_hd__o21bai_2 _5004_ (.A1(_0764_),
    .A2(_0771_),
    .B1_N(_0772_),
    .Y(_0773_));
 sky130_fd_sc_hd__xnor2_1 _5005_ (.A(_0764_),
    .B(_0771_),
    .Y(_0774_));
 sky130_fd_sc_hd__nand2_1 _5006_ (.A(_0774_),
    .B(_0772_),
    .Y(_0775_));
 sky130_fd_sc_hd__o21ai_2 _5007_ (.A1(_0770_),
    .A2(_0773_),
    .B1(_0775_),
    .Y(_0776_));
 sky130_fd_sc_hd__nand2_1 _5008_ (.A(_0709_),
    .B(_0748_),
    .Y(_0777_));
 sky130_fd_sc_hd__nor2_1 _5009_ (.A(_0710_),
    .B(_0749_),
    .Y(_0778_));
 sky130_fd_sc_hd__a22oi_2 _5010_ (.A1(_0747_),
    .A2(_0777_),
    .B1(_0655_),
    .B2(_0778_),
    .Y(_0779_));
 sky130_fd_sc_hd__xor2_1 _5011_ (.A(_0776_),
    .B(_0779_),
    .X(_0080_));
 sky130_fd_sc_hd__o22ai_1 _5012_ (.A1(_0770_),
    .A2(_0773_),
    .B1(_0776_),
    .B2(_0779_),
    .Y(_0780_));
 sky130_fd_sc_hd__mux2_1 _5013_ (.A0(_0762_),
    .A1(_0761_),
    .S(_0739_),
    .X(_0781_));
 sky130_fd_sc_hd__mux2_1 _5014_ (.A0(_0757_),
    .A1(_0758_),
    .S(_0664_),
    .X(_0782_));
 sky130_fd_sc_hd__xnor2_1 _5015_ (.A(_0764_),
    .B(_0754_),
    .Y(_0783_));
 sky130_fd_sc_hd__xor2_1 _5016_ (.A(_0782_),
    .B(_0783_),
    .X(_0784_));
 sky130_fd_sc_hd__xnor2_1 _5017_ (.A(_0781_),
    .B(_0784_),
    .Y(_0785_));
 sky130_fd_sc_hd__a21oi_1 _5018_ (.A1(_0769_),
    .A2(_0764_),
    .B1(_0768_),
    .Y(_0786_));
 sky130_fd_sc_hd__xnor2_1 _5019_ (.A(_0785_),
    .B(_0786_),
    .Y(_0787_));
 sky130_fd_sc_hd__nand2_1 _5020_ (.A(_0780_),
    .B(_0787_),
    .Y(_0788_));
 sky130_fd_sc_hd__xor2_1 _5021_ (.A(_0785_),
    .B(_0786_),
    .X(_0789_));
 sky130_fd_sc_hd__a21o_1 _5022_ (.A1(_0764_),
    .A2(_0771_),
    .B1(_0773_),
    .X(_0790_));
 sky130_fd_sc_hd__o211ai_1 _5023_ (.A1(_0776_),
    .A2(_0779_),
    .B1(_0789_),
    .C1(_0790_),
    .Y(_0791_));
 sky130_fd_sc_hd__nand2_1 _5024_ (.A(_0788_),
    .B(_0791_),
    .Y(_0081_));
 sky130_fd_sc_hd__a21bo_1 _5025_ (.A1(_0421_),
    .A2(_0420_),
    .B1_N(_0439_),
    .X(_0792_));
 sky130_fd_sc_hd__xor2_1 _5026_ (.A(_0436_),
    .B(_0792_),
    .X(_0067_));
 sky130_fd_sc_hd__and2_1 _5027_ (.A(\mixer_i.nco_valid ),
    .B(net531),
    .X(_0793_));
 sky130_fd_sc_hd__clkbuf_1 _5028_ (.A(net532),
    .X(_0024_));
 sky130_fd_sc_hd__inv_2 _5029_ (.A(net420),
    .Y(_0794_));
 sky130_fd_sc_hd__buf_2 _5030_ (.A(_0794_),
    .X(_0795_));
 sky130_fd_sc_hd__nand2_2 _5031_ (.A(_0795_),
    .B(net413),
    .Y(_0796_));
 sky130_fd_sc_hd__inv_2 _5032_ (.A(net461),
    .Y(_0797_));
 sky130_fd_sc_hd__inv_2 _5033_ (.A(net454),
    .Y(_0798_));
 sky130_fd_sc_hd__nor2_1 _5034_ (.A(_0797_),
    .B(_0798_),
    .Y(_0799_));
 sky130_fd_sc_hd__clkbuf_4 _5035_ (.A(_0799_),
    .X(_0800_));
 sky130_fd_sc_hd__o21ai_1 _5036_ (.A1(net459),
    .A2(net442),
    .B1(net427),
    .Y(_0801_));
 sky130_fd_sc_hd__clkbuf_4 _5037_ (.A(_0801_),
    .X(_0802_));
 sky130_fd_sc_hd__buf_4 _5038_ (.A(_0797_),
    .X(_0803_));
 sky130_fd_sc_hd__nand2_4 _5039_ (.A(_0803_),
    .B(_0798_),
    .Y(_0804_));
 sky130_fd_sc_hd__nand2_1 _5040_ (.A(net459),
    .B(net452),
    .Y(_0805_));
 sky130_fd_sc_hd__buf_2 _5041_ (.A(_0805_),
    .X(_0806_));
 sky130_fd_sc_hd__and3_1 _5042_ (.A(_0804_),
    .B(net443),
    .C(_0806_),
    .X(_0807_));
 sky130_fd_sc_hd__o32a_1 _5043_ (.A1(net426),
    .A2(net443),
    .A3(_0800_),
    .B1(_0802_),
    .B2(_0807_),
    .X(_0808_));
 sky130_fd_sc_hd__nor2_4 _5044_ (.A(net446),
    .B(_0803_),
    .Y(_0809_));
 sky130_fd_sc_hd__clkbuf_4 _5045_ (.A(_0803_),
    .X(_0810_));
 sky130_fd_sc_hd__a31o_1 _5046_ (.A1(_0810_),
    .A2(net452),
    .A3(net443),
    .B1(_0794_),
    .X(_0811_));
 sky130_fd_sc_hd__clkbuf_4 _5047_ (.A(_0810_),
    .X(_0812_));
 sky130_fd_sc_hd__clkbuf_4 _5048_ (.A(_0798_),
    .X(_0813_));
 sky130_fd_sc_hd__clkbuf_4 _5049_ (.A(_0813_),
    .X(_0814_));
 sky130_fd_sc_hd__buf_4 _5050_ (.A(_0814_),
    .X(_0815_));
 sky130_fd_sc_hd__inv_2 _5051_ (.A(net443),
    .Y(_0816_));
 sky130_fd_sc_hd__buf_2 _5052_ (.A(_0816_),
    .X(_0817_));
 sky130_fd_sc_hd__clkbuf_4 _5053_ (.A(_0817_),
    .X(_0818_));
 sky130_fd_sc_hd__clkbuf_4 _5054_ (.A(_0818_),
    .X(_0819_));
 sky130_fd_sc_hd__o21ai_2 _5055_ (.A1(_0810_),
    .A2(_0814_),
    .B1(net425),
    .Y(_0820_));
 sky130_fd_sc_hd__buf_4 _5056_ (.A(_0795_),
    .X(_0821_));
 sky130_fd_sc_hd__a311o_1 _5057_ (.A1(_0812_),
    .A2(_0815_),
    .A3(_0819_),
    .B1(_0820_),
    .C1(_0821_),
    .X(_0822_));
 sky130_fd_sc_hd__inv_2 _5058_ (.A(net426),
    .Y(_0823_));
 sky130_fd_sc_hd__nor2_4 _5059_ (.A(net414),
    .B(_0823_),
    .Y(_0824_));
 sky130_fd_sc_hd__a21oi_1 _5060_ (.A1(net459),
    .A2(net452),
    .B1(_0816_),
    .Y(_0825_));
 sky130_fd_sc_hd__a21o_1 _5061_ (.A1(net452),
    .A2(_0809_),
    .B1(_0825_),
    .X(_0826_));
 sky130_fd_sc_hd__nor2_4 _5062_ (.A(net459),
    .B(net442),
    .Y(_0827_));
 sky130_fd_sc_hd__nor2_2 _5063_ (.A(_0813_),
    .B(_0817_),
    .Y(_0828_));
 sky130_fd_sc_hd__nor2_4 _5064_ (.A(net453),
    .B(net447),
    .Y(_0829_));
 sky130_fd_sc_hd__or4_1 _5065_ (.A(net420),
    .B(_0827_),
    .C(_0828_),
    .D(_0829_),
    .X(_0830_));
 sky130_fd_sc_hd__a221o_1 _5066_ (.A1(_0824_),
    .A2(_0826_),
    .B1(_0830_),
    .B2(_0823_),
    .C1(net408),
    .X(_0831_));
 sky130_fd_sc_hd__o311a_1 _5067_ (.A1(net426),
    .A2(_0809_),
    .A3(_0811_),
    .B1(_0822_),
    .C1(_0831_),
    .X(_0832_));
 sky130_fd_sc_hd__o21ai_2 _5068_ (.A1(_0796_),
    .A2(_0808_),
    .B1(_0832_),
    .Y(_0833_));
 sky130_fd_sc_hd__inv_2 _5069_ (.A(net410),
    .Y(_0834_));
 sky130_fd_sc_hd__clkbuf_4 _5070_ (.A(_0834_),
    .X(_0835_));
 sky130_fd_sc_hd__buf_2 _5071_ (.A(_0835_),
    .X(_0836_));
 sky130_fd_sc_hd__nor2_2 _5072_ (.A(net431),
    .B(net458),
    .Y(_0837_));
 sky130_fd_sc_hd__nand2_4 _5073_ (.A(_0803_),
    .B(_0816_),
    .Y(_0838_));
 sky130_fd_sc_hd__nand2_2 _5074_ (.A(net458),
    .B(net444),
    .Y(_0839_));
 sky130_fd_sc_hd__and3_2 _5075_ (.A(_0838_),
    .B(_0839_),
    .C(net428),
    .X(_0840_));
 sky130_fd_sc_hd__or2_1 _5076_ (.A(net430),
    .B(_0814_),
    .X(_0841_));
 sky130_fd_sc_hd__or4b_1 _5077_ (.A(net417),
    .B(_0837_),
    .C(_0840_),
    .D_N(_0841_),
    .X(_0842_));
 sky130_fd_sc_hd__nand2_1 _5078_ (.A(net452),
    .B(net442),
    .Y(_0843_));
 sky130_fd_sc_hd__clkbuf_4 _5079_ (.A(_0843_),
    .X(_0844_));
 sky130_fd_sc_hd__buf_2 _5080_ (.A(_0844_),
    .X(_0845_));
 sky130_fd_sc_hd__o221ai_1 _5081_ (.A1(net437),
    .A2(net455),
    .B1(_0845_),
    .B2(_0837_),
    .C1(net422),
    .Y(_0846_));
 sky130_fd_sc_hd__clkbuf_4 _5082_ (.A(_0804_),
    .X(_0847_));
 sky130_fd_sc_hd__buf_2 _5083_ (.A(_0839_),
    .X(_0848_));
 sky130_fd_sc_hd__nand2_1 _5084_ (.A(_0838_),
    .B(_0848_),
    .Y(_0849_));
 sky130_fd_sc_hd__a21oi_1 _5085_ (.A1(_0814_),
    .A2(_0818_),
    .B1(net436),
    .Y(_0850_));
 sky130_fd_sc_hd__a31o_1 _5086_ (.A1(_0850_),
    .A2(net420),
    .A3(_0844_),
    .B1(_0834_),
    .X(_0851_));
 sky130_fd_sc_hd__nor2_4 _5087_ (.A(net460),
    .B(_0813_),
    .Y(_0852_));
 sky130_fd_sc_hd__clkbuf_4 _5088_ (.A(_0817_),
    .X(_0853_));
 sky130_fd_sc_hd__and3_1 _5089_ (.A(_0813_),
    .B(_0853_),
    .C(net460),
    .X(_0854_));
 sky130_fd_sc_hd__and3_1 _5090_ (.A(net462),
    .B(net456),
    .C(net446),
    .X(_0855_));
 sky130_fd_sc_hd__o311a_2 _5091_ (.A1(_0852_),
    .A2(_0854_),
    .A3(_0855_),
    .B1(net434),
    .C1(net421),
    .X(_0856_));
 sky130_fd_sc_hd__a311oi_1 _5092_ (.A1(_0824_),
    .A2(_0847_),
    .A3(_0849_),
    .B1(_0851_),
    .C1(_0856_),
    .Y(_0857_));
 sky130_fd_sc_hd__a31o_1 _5093_ (.A1(_0836_),
    .A2(_0842_),
    .A3(_0846_),
    .B1(_0857_),
    .X(_0858_));
 sky130_fd_sc_hd__inv_2 _5094_ (.A(net402),
    .Y(_0859_));
 sky130_fd_sc_hd__buf_2 _5095_ (.A(_0859_),
    .X(_0860_));
 sky130_fd_sc_hd__buf_2 _5096_ (.A(_0860_),
    .X(_0861_));
 sky130_fd_sc_hd__mux2_1 _5097_ (.A0(_0833_),
    .A1(_0858_),
    .S(_0861_),
    .X(_0862_));
 sky130_fd_sc_hd__clkbuf_1 _5098_ (.A(_0862_),
    .X(_0000_));
 sky130_fd_sc_hd__clkbuf_4 _5099_ (.A(_0794_),
    .X(_0863_));
 sky130_fd_sc_hd__buf_4 _5100_ (.A(_0863_),
    .X(_0864_));
 sky130_fd_sc_hd__nand2_2 _5101_ (.A(_0817_),
    .B(net461),
    .Y(_0865_));
 sky130_fd_sc_hd__a21oi_4 _5102_ (.A1(_0803_),
    .A2(net446),
    .B1(net454),
    .Y(_0866_));
 sky130_fd_sc_hd__and2b_1 _5103_ (.A_N(net425),
    .B(_0826_),
    .X(_0867_));
 sky130_fd_sc_hd__a31o_1 _5104_ (.A1(net436),
    .A2(_0865_),
    .A3(_0866_),
    .B1(_0867_),
    .X(_0868_));
 sky130_fd_sc_hd__nand2_2 _5105_ (.A(net426),
    .B(net452),
    .Y(_0869_));
 sky130_fd_sc_hd__a22o_2 _5106_ (.A1(net443),
    .A2(_0805_),
    .B1(_0801_),
    .B2(_0869_),
    .X(_0870_));
 sky130_fd_sc_hd__a31o_1 _5107_ (.A1(net460),
    .A2(net453),
    .A3(_0818_),
    .B1(_0870_),
    .X(_0871_));
 sky130_fd_sc_hd__o21a_1 _5108_ (.A1(net435),
    .A2(net460),
    .B1(_0795_),
    .X(_0872_));
 sky130_fd_sc_hd__a2bb2o_1 _5109_ (.A1_N(_0864_),
    .A2_N(_0868_),
    .B1(_0871_),
    .B2(_0872_),
    .X(_0873_));
 sky130_fd_sc_hd__or3_1 _5110_ (.A(net433),
    .B(_0810_),
    .C(_0829_),
    .X(_0874_));
 sky130_fd_sc_hd__clkbuf_4 _5111_ (.A(_0814_),
    .X(_0875_));
 sky130_fd_sc_hd__o21ai_1 _5112_ (.A1(_0875_),
    .A2(_0848_),
    .B1(net437),
    .Y(_0876_));
 sky130_fd_sc_hd__and4_1 _5113_ (.A(_0874_),
    .B(net422),
    .C(net412),
    .D(_0876_),
    .X(_0877_));
 sky130_fd_sc_hd__nand2_2 _5114_ (.A(_0810_),
    .B(net453),
    .Y(_0878_));
 sky130_fd_sc_hd__a32o_1 _5115_ (.A1(net439),
    .A2(net455),
    .A3(net448),
    .B1(_0878_),
    .B2(_0802_),
    .X(_0879_));
 sky130_fd_sc_hd__and3_1 _5116_ (.A(_0879_),
    .B(net413),
    .C(_0821_),
    .X(_0880_));
 sky130_fd_sc_hd__a211o_1 _5117_ (.A1(_0836_),
    .A2(_0873_),
    .B1(_0877_),
    .C1(_0880_),
    .X(_0881_));
 sky130_fd_sc_hd__o22a_1 _5118_ (.A1(_0813_),
    .A2(_0838_),
    .B1(_0817_),
    .B2(_0852_),
    .X(_0882_));
 sky130_fd_sc_hd__a31o_1 _5119_ (.A1(_0812_),
    .A2(net455),
    .A3(_0819_),
    .B1(_0876_),
    .X(_0883_));
 sky130_fd_sc_hd__o211a_1 _5120_ (.A1(net433),
    .A2(_0882_),
    .B1(_0883_),
    .C1(net420),
    .X(_0884_));
 sky130_fd_sc_hd__nor2_4 _5121_ (.A(net461),
    .B(_0817_),
    .Y(_0885_));
 sky130_fd_sc_hd__buf_2 _5122_ (.A(_0885_),
    .X(_0886_));
 sky130_fd_sc_hd__a31o_1 _5123_ (.A1(_0886_),
    .A2(_0795_),
    .A3(net438),
    .B1(net412),
    .X(_0887_));
 sky130_fd_sc_hd__a31o_1 _5124_ (.A1(_0821_),
    .A2(_0815_),
    .A3(_0849_),
    .B1(_0887_),
    .X(_0888_));
 sky130_fd_sc_hd__a21oi_4 _5125_ (.A1(_0818_),
    .A2(net463),
    .B1(net433),
    .Y(_0889_));
 sky130_fd_sc_hd__nor2_1 _5126_ (.A(net461),
    .B(net454),
    .Y(_0890_));
 sky130_fd_sc_hd__nor2_2 _5127_ (.A(_0799_),
    .B(_0890_),
    .Y(_0891_));
 sky130_fd_sc_hd__nand2_4 _5128_ (.A(net407),
    .B(net414),
    .Y(_0892_));
 sky130_fd_sc_hd__and3_4 _5129_ (.A(_0803_),
    .B(_0813_),
    .C(_0817_),
    .X(_0893_));
 sky130_fd_sc_hd__a221o_1 _5130_ (.A1(_0853_),
    .A2(net453),
    .B1(_0866_),
    .B2(_0865_),
    .C1(_0852_),
    .X(_0894_));
 sky130_fd_sc_hd__o21a_1 _5131_ (.A1(net435),
    .A2(_0893_),
    .B1(_0894_),
    .X(_0895_));
 sky130_fd_sc_hd__o32a_1 _5132_ (.A1(_0796_),
    .A2(_0889_),
    .A3(_0891_),
    .B1(_0892_),
    .B2(_0895_),
    .X(_0896_));
 sky130_fd_sc_hd__o21ai_2 _5133_ (.A1(_0884_),
    .A2(_0888_),
    .B1(_0896_),
    .Y(_0897_));
 sky130_fd_sc_hd__nand2_4 _5134_ (.A(_0805_),
    .B(_0804_),
    .Y(_0898_));
 sky130_fd_sc_hd__a32o_1 _5135_ (.A1(_0845_),
    .A2(_0848_),
    .A3(_0850_),
    .B1(_0898_),
    .B2(_0819_),
    .X(_0899_));
 sky130_fd_sc_hd__o211a_1 _5136_ (.A1(_0814_),
    .A2(_0838_),
    .B1(_0839_),
    .C1(net425),
    .X(_0900_));
 sky130_fd_sc_hd__clkbuf_4 _5137_ (.A(_0829_),
    .X(_0901_));
 sky130_fd_sc_hd__a211o_1 _5138_ (.A1(net442),
    .A2(_0852_),
    .B1(_0901_),
    .C1(net427),
    .X(_0902_));
 sky130_fd_sc_hd__and4b_1 _5139_ (.A_N(_0900_),
    .B(net408),
    .C(_0821_),
    .D(_0902_),
    .X(_0903_));
 sky130_fd_sc_hd__clkbuf_4 _5140_ (.A(_0869_),
    .X(_0904_));
 sky130_fd_sc_hd__a31o_1 _5141_ (.A1(_0894_),
    .A2(_0802_),
    .A3(_0904_),
    .B1(net421),
    .X(_0905_));
 sky130_fd_sc_hd__nor3_1 _5142_ (.A(net426),
    .B(net459),
    .C(net442),
    .Y(_0906_));
 sky130_fd_sc_hd__or4_1 _5143_ (.A(_0863_),
    .B(net452),
    .C(_0840_),
    .D(_0906_),
    .X(_0907_));
 sky130_fd_sc_hd__and3_1 _5144_ (.A(_0835_),
    .B(_0905_),
    .C(_0907_),
    .X(_0908_));
 sky130_fd_sc_hd__a311oi_4 _5145_ (.A1(net408),
    .A2(net420),
    .A3(_0899_),
    .B1(_0903_),
    .C1(_0908_),
    .Y(_0909_));
 sky130_fd_sc_hd__o21ai_1 _5146_ (.A1(net462),
    .A2(_0815_),
    .B1(net438),
    .Y(_0910_));
 sky130_fd_sc_hd__o311a_1 _5147_ (.A1(net438),
    .A2(net448),
    .A3(_0800_),
    .B1(_0910_),
    .C1(net423),
    .X(_0911_));
 sky130_fd_sc_hd__or2_4 _5148_ (.A(net434),
    .B(net456),
    .X(_0912_));
 sky130_fd_sc_hd__o21ai_1 _5149_ (.A1(net448),
    .A2(_0812_),
    .B1(net439),
    .Y(_0913_));
 sky130_fd_sc_hd__o221a_1 _5150_ (.A1(net448),
    .A2(_0912_),
    .B1(_0913_),
    .B2(_0866_),
    .C1(_0821_),
    .X(_0914_));
 sky130_fd_sc_hd__clkbuf_4 _5151_ (.A(_0828_),
    .X(_0915_));
 sky130_fd_sc_hd__a21o_2 _5152_ (.A1(net434),
    .A2(net461),
    .B1(_0794_),
    .X(_0916_));
 sky130_fd_sc_hd__a21oi_1 _5153_ (.A1(_0866_),
    .A2(net439),
    .B1(_0916_),
    .Y(_0917_));
 sky130_fd_sc_hd__o31a_1 _5154_ (.A1(net439),
    .A2(_0915_),
    .A3(_0854_),
    .B1(_0917_),
    .X(_0918_));
 sky130_fd_sc_hd__o41ai_2 _5155_ (.A1(net423),
    .A2(_0915_),
    .A3(_0889_),
    .A4(_0854_),
    .B1(net412),
    .Y(_0919_));
 sky130_fd_sc_hd__o32ai_2 _5156_ (.A1(net413),
    .A2(_0911_),
    .A3(_0914_),
    .B1(_0918_),
    .B2(_0919_),
    .Y(_0920_));
 sky130_fd_sc_hd__inv_2 _5157_ (.A(net399),
    .Y(_0921_));
 sky130_fd_sc_hd__buf_2 _5158_ (.A(_0921_),
    .X(_0922_));
 sky130_fd_sc_hd__mux4_1 _5159_ (.A0(_0881_),
    .A1(_0897_),
    .A2(_0909_),
    .A3(_0920_),
    .S0(_0861_),
    .S1(_0922_),
    .X(_0923_));
 sky130_fd_sc_hd__clkbuf_1 _5160_ (.A(_0923_),
    .X(_0003_));
 sky130_fd_sc_hd__nor2_1 _5161_ (.A(_0859_),
    .B(_0921_),
    .Y(_0924_));
 sky130_fd_sc_hd__clkbuf_2 _5162_ (.A(_0924_),
    .X(_0925_));
 sky130_fd_sc_hd__and4_1 _5163_ (.A(_0864_),
    .B(_0912_),
    .C(_0904_),
    .D(_0802_),
    .X(_0926_));
 sky130_fd_sc_hd__buf_2 _5164_ (.A(_0890_),
    .X(_0927_));
 sky130_fd_sc_hd__or3_1 _5165_ (.A(_0828_),
    .B(_0829_),
    .C(_0927_),
    .X(_0928_));
 sky130_fd_sc_hd__a31o_1 _5166_ (.A1(_0928_),
    .A2(net423),
    .A3(_0910_),
    .B1(net412),
    .X(_0929_));
 sky130_fd_sc_hd__a21oi_1 _5167_ (.A1(net455),
    .A2(net448),
    .B1(net438),
    .Y(_0930_));
 sky130_fd_sc_hd__o32a_1 _5168_ (.A1(net438),
    .A2(_0800_),
    .A3(_0927_),
    .B1(_0886_),
    .B2(_0915_),
    .X(_0931_));
 sky130_fd_sc_hd__a211o_1 _5169_ (.A1(_0930_),
    .A2(_0891_),
    .B1(_0892_),
    .C1(_0931_),
    .X(_0932_));
 sky130_fd_sc_hd__or3_2 _5170_ (.A(net455),
    .B(net446),
    .C(_0810_),
    .X(_0933_));
 sky130_fd_sc_hd__o221a_1 _5171_ (.A1(_0875_),
    .A2(_0848_),
    .B1(_0869_),
    .B2(_0819_),
    .C1(_0933_),
    .X(_0934_));
 sky130_fd_sc_hd__a311o_1 _5172_ (.A1(net433),
    .A2(net446),
    .A3(_0800_),
    .B1(_0796_),
    .C1(_0934_),
    .X(_0935_));
 sky130_fd_sc_hd__o211a_1 _5173_ (.A1(_0926_),
    .A2(_0929_),
    .B1(_0932_),
    .C1(_0935_),
    .X(_0936_));
 sky130_fd_sc_hd__o21ai_2 _5174_ (.A1(net435),
    .A2(_0815_),
    .B1(_0871_),
    .Y(_0937_));
 sky130_fd_sc_hd__o221a_1 _5175_ (.A1(net414),
    .A2(_0808_),
    .B1(_0906_),
    .B2(_0937_),
    .C1(_0835_),
    .X(_0938_));
 sky130_fd_sc_hd__nor2_1 _5176_ (.A(net415),
    .B(_0834_),
    .Y(_0939_));
 sky130_fd_sc_hd__a211o_1 _5177_ (.A1(net451),
    .A2(_0819_),
    .B1(_0802_),
    .C1(_0852_),
    .X(_0940_));
 sky130_fd_sc_hd__o311a_1 _5178_ (.A1(net430),
    .A2(net458),
    .A3(net445),
    .B1(_0939_),
    .C1(_0940_),
    .X(_0941_));
 sky130_fd_sc_hd__nor2_2 _5179_ (.A(net426),
    .B(_0803_),
    .Y(_0942_));
 sky130_fd_sc_hd__o311a_1 _5180_ (.A1(net457),
    .A2(_0886_),
    .A3(_0942_),
    .B1(net417),
    .C1(net411),
    .X(_0943_));
 sky130_fd_sc_hd__or3_1 _5181_ (.A(_0938_),
    .B(_0941_),
    .C(_0943_),
    .X(_0944_));
 sky130_fd_sc_hd__and3_1 _5182_ (.A(_0861_),
    .B(_0944_),
    .C(net400),
    .X(_0945_));
 sky130_fd_sc_hd__nand2_2 _5183_ (.A(_0921_),
    .B(net404),
    .Y(_0946_));
 sky130_fd_sc_hd__a22o_1 _5184_ (.A1(_0898_),
    .A2(net437),
    .B1(_0933_),
    .B2(_0930_),
    .X(_0947_));
 sky130_fd_sc_hd__o21a_1 _5185_ (.A1(_0915_),
    .A2(_0901_),
    .B1(_0837_),
    .X(_0948_));
 sky130_fd_sc_hd__a311oi_1 _5186_ (.A1(net440),
    .A2(_0891_),
    .A3(_0845_),
    .B1(_0892_),
    .C1(_0948_),
    .Y(_0949_));
 sky130_fd_sc_hd__a221o_1 _5187_ (.A1(net451),
    .A2(_0812_),
    .B1(_0841_),
    .B2(_0838_),
    .C1(net417),
    .X(_0950_));
 sky130_fd_sc_hd__a221o_1 _5188_ (.A1(net440),
    .A2(_0845_),
    .B1(_0891_),
    .B2(_0889_),
    .C1(_0916_),
    .X(_0951_));
 sky130_fd_sc_hd__a21oi_1 _5189_ (.A1(_0950_),
    .A2(_0951_),
    .B1(net410),
    .Y(_0952_));
 sky130_fd_sc_hd__a211o_1 _5190_ (.A1(_0939_),
    .A2(_0947_),
    .B1(_0949_),
    .C1(_0952_),
    .X(_0953_));
 sky130_fd_sc_hd__nand2_4 _5191_ (.A(_0813_),
    .B(_0853_),
    .Y(_0954_));
 sky130_fd_sc_hd__o22a_1 _5192_ (.A1(_0812_),
    .A2(_0954_),
    .B1(_0848_),
    .B2(_0875_),
    .X(_0955_));
 sky130_fd_sc_hd__or3_1 _5193_ (.A(net430),
    .B(net458),
    .C(net445),
    .X(_0956_));
 sky130_fd_sc_hd__a221o_1 _5194_ (.A1(_0955_),
    .A2(_0956_),
    .B1(_0942_),
    .B2(_0901_),
    .C1(_0864_),
    .X(_0957_));
 sky130_fd_sc_hd__o211a_1 _5195_ (.A1(_0839_),
    .A2(net457),
    .B1(_0838_),
    .C1(_0841_),
    .X(_0958_));
 sky130_fd_sc_hd__or3_1 _5196_ (.A(net419),
    .B(_0906_),
    .C(_0958_),
    .X(_0959_));
 sky130_fd_sc_hd__o21ai_1 _5197_ (.A1(net460),
    .A2(net453),
    .B1(net446),
    .Y(_0960_));
 sky130_fd_sc_hd__o221a_1 _5198_ (.A1(_0799_),
    .A2(_0960_),
    .B1(_0891_),
    .B2(net446),
    .C1(net436),
    .X(_0961_));
 sky130_fd_sc_hd__o211a_1 _5199_ (.A1(_0853_),
    .A2(_0804_),
    .B1(_0806_),
    .C1(net425),
    .X(_0962_));
 sky130_fd_sc_hd__a311o_1 _5200_ (.A1(_0812_),
    .A2(_0875_),
    .A3(_0819_),
    .B1(_0863_),
    .C1(_0962_),
    .X(_0963_));
 sky130_fd_sc_hd__o311a_1 _5201_ (.A1(net414),
    .A2(_0906_),
    .A3(_0961_),
    .B1(_0963_),
    .C1(net407),
    .X(_0964_));
 sky130_fd_sc_hd__a31o_1 _5202_ (.A1(_0836_),
    .A2(_0957_),
    .A3(_0959_),
    .B1(_0964_),
    .X(_0965_));
 sky130_fd_sc_hd__nor2_2 _5203_ (.A(net404),
    .B(net400),
    .Y(_0966_));
 sky130_fd_sc_hd__a2bb2o_1 _5204_ (.A1_N(_0946_),
    .A2_N(_0953_),
    .B1(_0965_),
    .B2(_0966_),
    .X(_0967_));
 sky130_fd_sc_hd__a211o_1 _5205_ (.A1(_0925_),
    .A2(_0936_),
    .B1(_0945_),
    .C1(_0967_),
    .X(_0004_));
 sky130_fd_sc_hd__nor2_1 _5206_ (.A(net427),
    .B(_0853_),
    .Y(_0968_));
 sky130_fd_sc_hd__nor2_2 _5207_ (.A(net425),
    .B(net442),
    .Y(_0969_));
 sky130_fd_sc_hd__o21a_1 _5208_ (.A1(_0812_),
    .A2(_0815_),
    .B1(_0969_),
    .X(_0970_));
 sky130_fd_sc_hd__a31o_1 _5209_ (.A1(net430),
    .A2(net458),
    .A3(_0845_),
    .B1(_0811_),
    .X(_0971_));
 sky130_fd_sc_hd__o32a_1 _5210_ (.A1(net415),
    .A2(_0968_),
    .A3(_0893_),
    .B1(_0970_),
    .B2(_0971_),
    .X(_0972_));
 sky130_fd_sc_hd__a22o_1 _5211_ (.A1(net437),
    .A2(net455),
    .B1(net448),
    .B2(net462),
    .X(_0973_));
 sky130_fd_sc_hd__and3_1 _5212_ (.A(_0973_),
    .B(net422),
    .C(_0912_),
    .X(_0974_));
 sky130_fd_sc_hd__a21oi_1 _5213_ (.A1(_0866_),
    .A2(net439),
    .B1(net422),
    .Y(_0975_));
 sky130_fd_sc_hd__a21o_1 _5214_ (.A1(_0866_),
    .A2(net440),
    .B1(net423),
    .X(_0976_));
 sky130_fd_sc_hd__a21oi_2 _5215_ (.A1(net437),
    .A2(net462),
    .B1(_0976_),
    .Y(_0977_));
 sky130_fd_sc_hd__a221o_1 _5216_ (.A1(net448),
    .A2(_0975_),
    .B1(_0977_),
    .B2(_0847_),
    .C1(_0834_),
    .X(_0978_));
 sky130_fd_sc_hd__o22a_1 _5217_ (.A1(net412),
    .A2(_0972_),
    .B1(_0974_),
    .B2(_0978_),
    .X(_0979_));
 sky130_fd_sc_hd__a21o_1 _5218_ (.A1(_0878_),
    .A2(net449),
    .B1(net438),
    .X(_0980_));
 sky130_fd_sc_hd__or3_1 _5219_ (.A(net462),
    .B(net455),
    .C(net448),
    .X(_0981_));
 sky130_fd_sc_hd__a21oi_1 _5220_ (.A1(_0981_),
    .A2(_0874_),
    .B1(_0795_),
    .Y(_0982_));
 sky130_fd_sc_hd__a21o_1 _5221_ (.A1(_0975_),
    .A2(_0980_),
    .B1(_0982_),
    .X(_0983_));
 sky130_fd_sc_hd__o32a_1 _5222_ (.A1(net438),
    .A2(_0901_),
    .A3(_0886_),
    .B1(_0913_),
    .B2(_0927_),
    .X(_0984_));
 sky130_fd_sc_hd__o2111ai_2 _5223_ (.A1(net437),
    .A2(_0893_),
    .B1(_0844_),
    .C1(net422),
    .D1(_0848_),
    .Y(_0985_));
 sky130_fd_sc_hd__o211a_1 _5224_ (.A1(net422),
    .A2(_0984_),
    .B1(_0985_),
    .C1(net412),
    .X(_0986_));
 sky130_fd_sc_hd__a21o_1 _5225_ (.A1(_0836_),
    .A2(_0983_),
    .B1(_0986_),
    .X(_0987_));
 sky130_fd_sc_hd__nor2_1 _5226_ (.A(net404),
    .B(_0921_),
    .Y(_0988_));
 sky130_fd_sc_hd__o22a_1 _5227_ (.A1(_0814_),
    .A2(net462),
    .B1(_0886_),
    .B2(_0828_),
    .X(_0989_));
 sky130_fd_sc_hd__a221o_1 _5228_ (.A1(_0824_),
    .A2(_0933_),
    .B1(_0989_),
    .B2(_0864_),
    .C1(_0982_),
    .X(_0990_));
 sky130_fd_sc_hd__o32a_1 _5229_ (.A1(net437),
    .A2(_0829_),
    .A3(_0885_),
    .B1(_0904_),
    .B2(_0809_),
    .X(_0991_));
 sky130_fd_sc_hd__o211a_1 _5230_ (.A1(net423),
    .A2(_0991_),
    .B1(_0985_),
    .C1(net412),
    .X(_0992_));
 sky130_fd_sc_hd__a21o_1 _5231_ (.A1(_0836_),
    .A2(_0990_),
    .B1(_0992_),
    .X(_0993_));
 sky130_fd_sc_hd__a31o_1 _5232_ (.A1(net428),
    .A2(_0815_),
    .A3(_0827_),
    .B1(_0968_),
    .X(_0994_));
 sky130_fd_sc_hd__o22ai_4 _5233_ (.A1(net415),
    .A2(_0994_),
    .B1(_0969_),
    .B2(_0971_),
    .Y(_0995_));
 sky130_fd_sc_hd__a211o_1 _5234_ (.A1(net458),
    .A2(net445),
    .B1(_0802_),
    .C1(_0852_),
    .X(_0996_));
 sky130_fd_sc_hd__and4b_1 _5235_ (.A_N(_0837_),
    .B(_0912_),
    .C(_0996_),
    .D(net423),
    .X(_0997_));
 sky130_fd_sc_hd__o2bb2a_1 _5236_ (.A1_N(_0836_),
    .A2_N(_0995_),
    .B1(_0997_),
    .B2(_0978_),
    .X(_0998_));
 sky130_fd_sc_hd__a22oi_1 _5237_ (.A1(_0988_),
    .A2(_0993_),
    .B1(_0998_),
    .B2(_0925_),
    .Y(_0999_));
 sky130_fd_sc_hd__o31a_1 _5238_ (.A1(net406),
    .A2(net401),
    .A3(_0987_),
    .B1(_0999_),
    .X(_1000_));
 sky130_fd_sc_hd__o21ai_1 _5239_ (.A1(_0946_),
    .A2(_0979_),
    .B1(net787),
    .Y(_0005_));
 sky130_fd_sc_hd__o311a_1 _5240_ (.A1(net451),
    .A2(_0809_),
    .A3(_0885_),
    .B1(_0806_),
    .C1(net430),
    .X(_1001_));
 sky130_fd_sc_hd__a21oi_1 _5241_ (.A1(_0844_),
    .A2(_0839_),
    .B1(net428),
    .Y(_1002_));
 sky130_fd_sc_hd__o21a_1 _5242_ (.A1(_1001_),
    .A2(_1002_),
    .B1(_0821_),
    .X(_1003_));
 sky130_fd_sc_hd__o31a_1 _5243_ (.A1(net431),
    .A2(_0901_),
    .A3(_0898_),
    .B1(net418),
    .X(_1004_));
 sky130_fd_sc_hd__a211o_1 _5244_ (.A1(_0865_),
    .A2(net437),
    .B1(net455),
    .C1(_0886_),
    .X(_1005_));
 sky130_fd_sc_hd__a21o_1 _5245_ (.A1(_0954_),
    .A2(_0837_),
    .B1(_0916_),
    .X(_1006_));
 sky130_fd_sc_hd__or4b_2 _5246_ (.A(net422),
    .B(net462),
    .C(_0818_),
    .D_N(_0912_),
    .X(_1007_));
 sky130_fd_sc_hd__o2111ai_4 _5247_ (.A1(net422),
    .A2(_1005_),
    .B1(net410),
    .C1(_1006_),
    .D1(_1007_),
    .Y(_1008_));
 sky130_fd_sc_hd__o31a_1 _5248_ (.A1(net410),
    .A2(_1003_),
    .A3(_1004_),
    .B1(_1008_),
    .X(_1009_));
 sky130_fd_sc_hd__and3_1 _5249_ (.A(net417),
    .B(_0942_),
    .C(_0845_),
    .X(_1010_));
 sky130_fd_sc_hd__o2111a_1 _5250_ (.A1(net445),
    .A2(_0875_),
    .B1(net430),
    .C1(net417),
    .D1(_0865_),
    .X(_1011_));
 sky130_fd_sc_hd__a311o_1 _5251_ (.A1(net451),
    .A2(_0824_),
    .A3(_0848_),
    .B1(_0834_),
    .C1(_1011_),
    .X(_1012_));
 sky130_fd_sc_hd__o32a_1 _5252_ (.A1(net430),
    .A2(_0809_),
    .A3(_0807_),
    .B1(_0886_),
    .B2(_0904_),
    .X(_1013_));
 sky130_fd_sc_hd__a21o_1 _5253_ (.A1(net417),
    .A2(_1013_),
    .B1(net410),
    .X(_1014_));
 sky130_fd_sc_hd__o31a_1 _5254_ (.A1(net431),
    .A2(net459),
    .A3(_0901_),
    .B1(_0977_),
    .X(_1015_));
 sky130_fd_sc_hd__o22a_1 _5255_ (.A1(_1010_),
    .A2(_1012_),
    .B1(_1014_),
    .B2(_1015_),
    .X(_1016_));
 sky130_fd_sc_hd__and3_1 _5256_ (.A(net417),
    .B(_0942_),
    .C(_0875_),
    .X(_1017_));
 sky130_fd_sc_hd__a31o_1 _5257_ (.A1(net417),
    .A2(net457),
    .A3(_0809_),
    .B1(_1017_),
    .X(_1018_));
 sky130_fd_sc_hd__o21a_1 _5258_ (.A1(net431),
    .A2(net458),
    .B1(_0977_),
    .X(_1019_));
 sky130_fd_sc_hd__o22a_1 _5259_ (.A1(_1012_),
    .A2(_1018_),
    .B1(_1014_),
    .B2(_1019_),
    .X(_1020_));
 sky130_fd_sc_hd__nor2_1 _5260_ (.A(net430),
    .B(_0845_),
    .Y(_1021_));
 sky130_fd_sc_hd__o21a_1 _5261_ (.A1(_1001_),
    .A2(_1021_),
    .B1(_0864_),
    .X(_1022_));
 sky130_fd_sc_hd__o31a_1 _5262_ (.A1(net410),
    .A2(_1004_),
    .A3(_1022_),
    .B1(_1008_),
    .X(_1023_));
 sky130_fd_sc_hd__nand2_1 _5263_ (.A(_0860_),
    .B(_0921_),
    .Y(_1024_));
 sky130_fd_sc_hd__o2bb2a_1 _5264_ (.A1_N(_0925_),
    .A2_N(_1020_),
    .B1(_1023_),
    .B2(_1024_),
    .X(_1025_));
 sky130_fd_sc_hd__o21ai_1 _5265_ (.A1(_0946_),
    .A2(_1016_),
    .B1(_1025_),
    .Y(_1026_));
 sky130_fd_sc_hd__a31o_1 _5266_ (.A1(_0861_),
    .A2(net400),
    .A3(_1009_),
    .B1(_1026_),
    .X(_0006_));
 sky130_fd_sc_hd__or2_1 _5267_ (.A(_0925_),
    .B(_0966_),
    .X(_1027_));
 sky130_fd_sc_hd__nor2_1 _5268_ (.A(_0924_),
    .B(_0966_),
    .Y(_1028_));
 sky130_fd_sc_hd__o41a_1 _5269_ (.A1(net416),
    .A2(net429),
    .A3(net444),
    .A4(_0847_),
    .B1(_1028_),
    .X(_1029_));
 sky130_fd_sc_hd__a311oi_2 _5270_ (.A1(_0843_),
    .A2(_0954_),
    .A3(_0804_),
    .B1(_0893_),
    .C1(net427),
    .Y(_1030_));
 sky130_fd_sc_hd__o221a_1 _5271_ (.A1(net414),
    .A2(_0962_),
    .B1(_0916_),
    .B2(_1030_),
    .C1(_0835_),
    .X(_1031_));
 sky130_fd_sc_hd__o2111a_1 _5272_ (.A1(net428),
    .A2(_0898_),
    .B1(_0904_),
    .C1(net409),
    .D1(net415),
    .X(_1032_));
 sky130_fd_sc_hd__and2_2 _5273_ (.A(net425),
    .B(net442),
    .X(_1033_));
 sky130_fd_sc_hd__or4_1 _5274_ (.A(net451),
    .B(_0809_),
    .C(_1033_),
    .D(_0885_),
    .X(_1034_));
 sky130_fd_sc_hd__o22a_1 _5275_ (.A1(net444),
    .A2(_0806_),
    .B1(_0904_),
    .B2(_0827_),
    .X(_1035_));
 sky130_fd_sc_hd__and3_1 _5276_ (.A(_1034_),
    .B(_1035_),
    .C(_0939_),
    .X(_1036_));
 sky130_fd_sc_hd__and3_1 _5277_ (.A(_0912_),
    .B(net419),
    .C(net408),
    .X(_1037_));
 sky130_fd_sc_hd__o211a_1 _5278_ (.A1(_0942_),
    .A2(_0961_),
    .B1(net408),
    .C1(_0794_),
    .X(_1038_));
 sky130_fd_sc_hd__a31o_1 _5279_ (.A1(_0802_),
    .A2(_0904_),
    .A3(_1037_),
    .B1(_1038_),
    .X(_1039_));
 sky130_fd_sc_hd__a2111oi_2 _5280_ (.A1(_0853_),
    .A2(net436),
    .B1(_0927_),
    .C1(_0800_),
    .D1(_0885_),
    .Y(_1040_));
 sky130_fd_sc_hd__a311oi_4 _5281_ (.A1(net436),
    .A2(_0818_),
    .A3(_0898_),
    .B1(_0863_),
    .C1(_1040_),
    .Y(_1041_));
 sky130_fd_sc_hd__o311a_1 _5282_ (.A1(net426),
    .A2(_0800_),
    .A3(_0927_),
    .B1(_0869_),
    .C1(_0794_),
    .X(_1042_));
 sky130_fd_sc_hd__o21a_1 _5283_ (.A1(_1041_),
    .A2(_1042_),
    .B1(_0834_),
    .X(_1043_));
 sky130_fd_sc_hd__or3_1 _5284_ (.A(_0859_),
    .B(_1039_),
    .C(_1043_),
    .X(_1044_));
 sky130_fd_sc_hd__o41a_1 _5285_ (.A1(net403),
    .A2(_1031_),
    .A3(_1032_),
    .A4(_1036_),
    .B1(_1044_),
    .X(_1045_));
 sky130_fd_sc_hd__mux2_1 _5286_ (.A0(_1027_),
    .A1(_1029_),
    .S(_1045_),
    .X(_1046_));
 sky130_fd_sc_hd__clkbuf_1 _5287_ (.A(_1046_),
    .X(_0007_));
 sky130_fd_sc_hd__or4_2 _5288_ (.A(net429),
    .B(net458),
    .C(net451),
    .D(net444),
    .X(_1047_));
 sky130_fd_sc_hd__o31a_1 _5289_ (.A1(net409),
    .A2(net416),
    .A3(_1047_),
    .B1(_1028_),
    .X(_1048_));
 sky130_fd_sc_hd__o311a_1 _5290_ (.A1(net433),
    .A2(_0800_),
    .A3(_0927_),
    .B1(_0870_),
    .C1(_0795_),
    .X(_1049_));
 sky130_fd_sc_hd__o21ai_1 _5291_ (.A1(net436),
    .A2(_0882_),
    .B1(_0863_),
    .Y(_1050_));
 sky130_fd_sc_hd__o21ai_1 _5292_ (.A1(net454),
    .A2(_0810_),
    .B1(net433),
    .Y(_1051_));
 sky130_fd_sc_hd__a32o_1 _5293_ (.A1(net433),
    .A2(net447),
    .A3(_0878_),
    .B1(_0882_),
    .B2(_1051_),
    .X(_1052_));
 sky130_fd_sc_hd__a2bb2o_1 _5294_ (.A1_N(_0961_),
    .A2_N(_1050_),
    .B1(_1052_),
    .B2(net420),
    .X(_1053_));
 sky130_fd_sc_hd__o22a_2 _5295_ (.A1(_0851_),
    .A2(_1049_),
    .B1(net413),
    .B2(_1053_),
    .X(_1054_));
 sky130_fd_sc_hd__a31o_1 _5296_ (.A1(_0806_),
    .A2(_0847_),
    .A3(_0889_),
    .B1(_0900_),
    .X(_1055_));
 sky130_fd_sc_hd__o211a_1 _5297_ (.A1(_0840_),
    .A2(_1030_),
    .B1(net407),
    .C1(net414),
    .X(_1056_));
 sky130_fd_sc_hd__o2111a_1 _5298_ (.A1(_0912_),
    .A2(_0885_),
    .B1(_0869_),
    .C1(_0844_),
    .D1(net414),
    .X(_1057_));
 sky130_fd_sc_hd__a311oi_4 _5299_ (.A1(_0864_),
    .A2(_0826_),
    .A3(net425),
    .B1(net407),
    .C1(_1057_),
    .Y(_1058_));
 sky130_fd_sc_hd__a311oi_4 _5300_ (.A1(net407),
    .A2(_0821_),
    .A3(_1055_),
    .B1(_1056_),
    .C1(_1058_),
    .Y(_1059_));
 sky130_fd_sc_hd__mux2_1 _5301_ (.A0(_1054_),
    .A1(_1059_),
    .S(_0860_),
    .X(_1060_));
 sky130_fd_sc_hd__mux2_1 _5302_ (.A0(_1027_),
    .A1(_1048_),
    .S(_1060_),
    .X(_1061_));
 sky130_fd_sc_hd__clkbuf_1 _5303_ (.A(_1061_),
    .X(_0008_));
 sky130_fd_sc_hd__a22o_1 _5304_ (.A1(_0825_),
    .A2(_0804_),
    .B1(_0898_),
    .B2(_0853_),
    .X(_1062_));
 sky130_fd_sc_hd__and4_1 _5305_ (.A(_0863_),
    .B(_1062_),
    .C(net426),
    .D(_0870_),
    .X(_1063_));
 sky130_fd_sc_hd__or4_1 _5306_ (.A(net436),
    .B(_0827_),
    .C(_0828_),
    .D(_0829_),
    .X(_1064_));
 sky130_fd_sc_hd__a22oi_1 _5307_ (.A1(_0824_),
    .A2(_1062_),
    .B1(_1064_),
    .B2(_0870_),
    .Y(_1065_));
 sky130_fd_sc_hd__a21o_1 _5308_ (.A1(_0969_),
    .A2(_0875_),
    .B1(_0863_),
    .X(_1066_));
 sky130_fd_sc_hd__o311ai_2 _5309_ (.A1(net414),
    .A2(_1033_),
    .A3(_0867_),
    .B1(_1066_),
    .C1(net407),
    .Y(_1067_));
 sky130_fd_sc_hd__o31a_2 _5310_ (.A1(net407),
    .A2(_1063_),
    .A3(_1065_),
    .B1(_1067_),
    .X(_1068_));
 sky130_fd_sc_hd__o311a_1 _5311_ (.A1(_0827_),
    .A2(_0915_),
    .A3(_0901_),
    .B1(net438),
    .C1(_0795_),
    .X(_1069_));
 sky130_fd_sc_hd__and4b_1 _5312_ (.A_N(net434),
    .B(_0960_),
    .C(_0954_),
    .D(_0794_),
    .X(_1070_));
 sky130_fd_sc_hd__a31o_1 _5313_ (.A1(net420),
    .A2(_0815_),
    .A3(_0889_),
    .B1(_1070_),
    .X(_1071_));
 sky130_fd_sc_hd__o21ai_1 _5314_ (.A1(_0828_),
    .A2(_0829_),
    .B1(net434),
    .Y(_1072_));
 sky130_fd_sc_hd__o311a_1 _5315_ (.A1(net433),
    .A2(_0818_),
    .A3(_0927_),
    .B1(net420),
    .C1(_1072_),
    .X(_1073_));
 sky130_fd_sc_hd__a311o_1 _5316_ (.A1(net462),
    .A2(_0824_),
    .A3(_0915_),
    .B1(_1073_),
    .C1(net412),
    .X(_1074_));
 sky130_fd_sc_hd__o41ai_4 _5317_ (.A1(_0835_),
    .A2(_0856_),
    .A3(_1069_),
    .A4(_1071_),
    .B1(_1074_),
    .Y(_1075_));
 sky130_fd_sc_hd__mux2_1 _5318_ (.A0(_1068_),
    .A1(_1075_),
    .S(_0860_),
    .X(_1076_));
 sky130_fd_sc_hd__mux2_1 _5319_ (.A0(_1029_),
    .A1(_1027_),
    .S(_1076_),
    .X(_1077_));
 sky130_fd_sc_hd__clkbuf_1 _5320_ (.A(_1077_),
    .X(_0009_));
 sky130_fd_sc_hd__o221a_1 _5321_ (.A1(net428),
    .A2(_0844_),
    .B1(_0820_),
    .B2(net444),
    .C1(_1047_),
    .X(_1078_));
 sky130_fd_sc_hd__a311o_1 _5322_ (.A1(net428),
    .A2(_0819_),
    .A3(_0806_),
    .B1(_1002_),
    .C1(net415),
    .X(_1079_));
 sky130_fd_sc_hd__a22o_1 _5323_ (.A1(net427),
    .A2(_0843_),
    .B1(_0968_),
    .B2(_0847_),
    .X(_1080_));
 sky130_fd_sc_hd__a21o_1 _5324_ (.A1(_1080_),
    .A2(net415),
    .B1(net407),
    .X(_1081_));
 sky130_fd_sc_hd__o211a_1 _5325_ (.A1(_0892_),
    .A2(_1078_),
    .B1(_1079_),
    .C1(_1081_),
    .X(_1082_));
 sky130_fd_sc_hd__a21o_1 _5326_ (.A1(_0969_),
    .A2(_0806_),
    .B1(_0834_),
    .X(_1083_));
 sky130_fd_sc_hd__o22a_1 _5327_ (.A1(net428),
    .A2(_0844_),
    .B1(net444),
    .B2(_0820_),
    .X(_1084_));
 sky130_fd_sc_hd__o21ai_2 _5328_ (.A1(net429),
    .A2(_0915_),
    .B1(net416),
    .Y(_1085_));
 sky130_fd_sc_hd__o2bb2a_1 _5329_ (.A1_N(_0864_),
    .A2_N(_1084_),
    .B1(_1085_),
    .B2(_1033_),
    .X(_1086_));
 sky130_fd_sc_hd__o32ai_2 _5330_ (.A1(net415),
    .A2(_1083_),
    .A3(_1033_),
    .B1(net409),
    .B2(_1086_),
    .Y(_1087_));
 sky130_fd_sc_hd__mux2_1 _5331_ (.A0(_1082_),
    .A1(_1087_),
    .S(net402),
    .X(_1088_));
 sky130_fd_sc_hd__a21bo_1 _5332_ (.A1(_1028_),
    .A2(_1047_),
    .B1_N(_1088_),
    .X(_1089_));
 sky130_fd_sc_hd__o31a_1 _5333_ (.A1(_0925_),
    .A2(_0966_),
    .A3(_1088_),
    .B1(_1089_),
    .X(_0010_));
 sky130_fd_sc_hd__a31o_1 _5334_ (.A1(_0838_),
    .A2(_0954_),
    .A3(net428),
    .B1(net415),
    .X(_1090_));
 sky130_fd_sc_hd__a2bb2o_1 _5335_ (.A1_N(_0835_),
    .A2_N(_0970_),
    .B1(_1085_),
    .B2(_1090_),
    .X(_1091_));
 sky130_fd_sc_hd__and3_1 _5336_ (.A(net429),
    .B(net451),
    .C(net444),
    .X(_1092_));
 sky130_fd_sc_hd__a2bb2o_1 _5337_ (.A1_N(net409),
    .A2_N(_1092_),
    .B1(_1085_),
    .B2(_1090_),
    .X(_1093_));
 sky130_fd_sc_hd__mux2_1 _5338_ (.A0(_1091_),
    .A1(_1093_),
    .S(_0860_),
    .X(_1094_));
 sky130_fd_sc_hd__mux2_1 _5339_ (.A0(_1048_),
    .A1(_1027_),
    .S(_1094_),
    .X(_1095_));
 sky130_fd_sc_hd__clkbuf_1 _5340_ (.A(_1095_),
    .X(_0011_));
 sky130_fd_sc_hd__and3_1 _5341_ (.A(_0859_),
    .B(_1090_),
    .C(net409),
    .X(_1096_));
 sky130_fd_sc_hd__a31o_1 _5342_ (.A1(net403),
    .A2(_0836_),
    .A3(_1085_),
    .B1(_1096_),
    .X(_1097_));
 sky130_fd_sc_hd__mux2_1 _5343_ (.A0(_1027_),
    .A1(_1029_),
    .S(_1097_),
    .X(_1098_));
 sky130_fd_sc_hd__clkbuf_1 _5344_ (.A(_1098_),
    .X(_0001_));
 sky130_fd_sc_hd__a21o_1 _5345_ (.A1(_0861_),
    .A2(net399),
    .B1(_1048_),
    .X(_0002_));
 sky130_fd_sc_hd__mux2_1 _5346_ (.A0(_0833_),
    .A1(_0858_),
    .S(net405),
    .X(_1099_));
 sky130_fd_sc_hd__clkbuf_1 _5347_ (.A(_1099_),
    .X(_0012_));
 sky130_fd_sc_hd__and3_1 _5348_ (.A(_0897_),
    .B(net401),
    .C(net406),
    .X(_1100_));
 sky130_fd_sc_hd__o32a_1 _5349_ (.A1(net966),
    .A2(_0911_),
    .A3(_0914_),
    .B1(_0918_),
    .B2(_0919_),
    .X(_1101_));
 sky130_fd_sc_hd__a2bb2o_1 _5350_ (.A1_N(_0946_),
    .A2_N(_1101_),
    .B1(_0966_),
    .B2(_0881_),
    .X(_1102_));
 sky130_fd_sc_hd__a211o_1 _5351_ (.A1(_0909_),
    .A2(_0988_),
    .B1(_1100_),
    .C1(_1102_),
    .X(_0015_));
 sky130_fd_sc_hd__and3_1 _5352_ (.A(_0936_),
    .B(_0921_),
    .C(_0861_),
    .X(_1103_));
 sky130_fd_sc_hd__and3_1 _5353_ (.A(_0965_),
    .B(net404),
    .C(_0922_),
    .X(_1104_));
 sky130_fd_sc_hd__nor3_1 _5354_ (.A(net404),
    .B(_0922_),
    .C(_0953_),
    .Y(_1105_));
 sky130_fd_sc_hd__a2111o_1 _5355_ (.A1(_0944_),
    .A2(_0925_),
    .B1(_1103_),
    .C1(_1104_),
    .D1(_1105_),
    .X(_0016_));
 sky130_fd_sc_hd__a22oi_1 _5356_ (.A1(_0925_),
    .A2(_0993_),
    .B1(_0998_),
    .B2(_0966_),
    .Y(_1106_));
 sky130_fd_sc_hd__o31a_1 _5357_ (.A1(_0861_),
    .A2(net401),
    .A3(_0987_),
    .B1(_1106_),
    .X(_1107_));
 sky130_fd_sc_hd__o31ai_1 _5358_ (.A1(net404),
    .A2(_0922_),
    .A3(_0979_),
    .B1(_1107_),
    .Y(_0017_));
 sky130_fd_sc_hd__nor3_1 _5359_ (.A(net404),
    .B(_0922_),
    .C(_1016_),
    .Y(_1108_));
 sky130_fd_sc_hd__a2bb2o_1 _5360_ (.A1_N(_0946_),
    .A2_N(_1023_),
    .B1(_1020_),
    .B2(_0966_),
    .X(_1109_));
 sky130_fd_sc_hd__a311o_1 _5361_ (.A1(net404),
    .A2(net400),
    .A3(_1009_),
    .B1(_1108_),
    .C1(_1109_),
    .X(_0018_));
 sky130_fd_sc_hd__or4_2 _5362_ (.A(net416),
    .B(net429),
    .C(net444),
    .D(_0847_),
    .X(_1110_));
 sky130_fd_sc_hd__o31a_1 _5363_ (.A1(net402),
    .A2(net410),
    .A3(_1110_),
    .B1(_0921_),
    .X(_1111_));
 sky130_fd_sc_hd__or4_1 _5364_ (.A(net425),
    .B(net451),
    .C(net442),
    .D(_1041_),
    .X(_1112_));
 sky130_fd_sc_hd__a211o_1 _5365_ (.A1(_1112_),
    .A2(_1043_),
    .B1(_1039_),
    .C1(net405),
    .X(_1113_));
 sky130_fd_sc_hd__o41ai_2 _5366_ (.A1(_0860_),
    .A2(_1031_),
    .A3(_1032_),
    .A4(_1036_),
    .B1(_1113_),
    .Y(_1114_));
 sky130_fd_sc_hd__mux2_1 _5367_ (.A0(net399),
    .A1(_1111_),
    .S(_1114_),
    .X(_1115_));
 sky130_fd_sc_hd__clkbuf_1 _5368_ (.A(_1115_),
    .X(_0019_));
 sky130_fd_sc_hd__o31a_1 _5369_ (.A1(net409),
    .A2(net416),
    .A3(_1047_),
    .B1(net399),
    .X(_1116_));
 sky130_fd_sc_hd__mux2_1 _5370_ (.A0(_1054_),
    .A1(_1059_),
    .S(net402),
    .X(_1117_));
 sky130_fd_sc_hd__mux2_1 _5371_ (.A0(_0922_),
    .A1(_1116_),
    .S(_1117_),
    .X(_1118_));
 sky130_fd_sc_hd__clkbuf_1 _5372_ (.A(_1118_),
    .X(_0020_));
 sky130_fd_sc_hd__mux2_1 _5373_ (.A0(_1068_),
    .A1(_1075_),
    .S(net403),
    .X(_1119_));
 sky130_fd_sc_hd__a21oi_1 _5374_ (.A1(net399),
    .A2(_1110_),
    .B1(_1119_),
    .Y(_1120_));
 sky130_fd_sc_hd__a21oi_1 _5375_ (.A1(net400),
    .A2(_1119_),
    .B1(_1120_),
    .Y(_0021_));
 sky130_fd_sc_hd__o31a_1 _5376_ (.A1(net429),
    .A2(net445),
    .A3(_0847_),
    .B1(_0860_),
    .X(_1121_));
 sky130_fd_sc_hd__a22o_1 _5377_ (.A1(_1087_),
    .A2(_1121_),
    .B1(_1082_),
    .B2(net402),
    .X(_1122_));
 sky130_fd_sc_hd__mux2_1 _5378_ (.A0(_1111_),
    .A1(net399),
    .S(_1122_),
    .X(_1123_));
 sky130_fd_sc_hd__clkbuf_1 _5379_ (.A(_1123_),
    .X(_0022_));
 sky130_fd_sc_hd__mux2_1 _5380_ (.A0(_1091_),
    .A1(_1093_),
    .S(net402),
    .X(_1124_));
 sky130_fd_sc_hd__mux2_1 _5381_ (.A0(_1116_),
    .A1(_0922_),
    .S(_1124_),
    .X(_1125_));
 sky130_fd_sc_hd__clkbuf_1 _5382_ (.A(_1125_),
    .X(_0023_));
 sky130_fd_sc_hd__and4_1 _5383_ (.A(_1085_),
    .B(_1110_),
    .C(_0835_),
    .D(_0859_),
    .X(_1126_));
 sky130_fd_sc_hd__a31o_1 _5384_ (.A1(net402),
    .A2(net409),
    .A3(_1090_),
    .B1(_1126_),
    .X(_1127_));
 sky130_fd_sc_hd__mux2_1 _5385_ (.A0(_1111_),
    .A1(net399),
    .S(_1127_),
    .X(_1128_));
 sky130_fd_sc_hd__clkbuf_1 _5386_ (.A(_1128_),
    .X(_0013_));
 sky130_fd_sc_hd__o31a_1 _5387_ (.A1(net402),
    .A2(net409),
    .A3(_1110_),
    .B1(net399),
    .X(_0014_));
 sky130_fd_sc_hd__clkinv_4 _5388_ (.A(net249),
    .Y(_1129_));
 sky130_fd_sc_hd__nor2_2 _5389_ (.A(_3125_),
    .B(_1129_),
    .Y(_0062_));
 sky130_fd_sc_hd__nor2_1 _5390_ (.A(net14),
    .B(net731),
    .Y(_1130_));
 sky130_fd_sc_hd__nand2_1 _5391_ (.A(net14),
    .B(\nco_inst.phase_accum[0] ),
    .Y(_1131_));
 sky130_fd_sc_hd__and2b_1 _5392_ (.A_N(_1130_),
    .B(net535),
    .X(_1132_));
 sky130_fd_sc_hd__clkbuf_1 _5393_ (.A(_1132_),
    .X(_0025_));
 sky130_fd_sc_hd__nor2_1 _5394_ (.A(net25),
    .B(\nco_inst.phase_accum[1] ),
    .Y(_1133_));
 sky130_fd_sc_hd__nand2_1 _5395_ (.A(net25),
    .B(\nco_inst.phase_accum[1] ),
    .Y(_1134_));
 sky130_fd_sc_hd__or2b_1 _5396_ (.A(_1133_),
    .B_N(_1134_),
    .X(_1135_));
 sky130_fd_sc_hd__xor2_1 _5397_ (.A(net535),
    .B(_1135_),
    .X(_0036_));
 sky130_fd_sc_hd__nor2_1 _5398_ (.A(net36),
    .B(\nco_inst.phase_accum[2] ),
    .Y(_1136_));
 sky130_fd_sc_hd__and2_1 _5399_ (.A(net36),
    .B(\nco_inst.phase_accum[2] ),
    .X(_1137_));
 sky130_fd_sc_hd__a22oi_2 _5400_ (.A1(net14),
    .A2(\nco_inst.phase_accum[0] ),
    .B1(net25),
    .B2(\nco_inst.phase_accum[1] ),
    .Y(_1138_));
 sky130_fd_sc_hd__or3_1 _5401_ (.A(_1133_),
    .B(_1137_),
    .C(_1138_),
    .X(_1139_));
 sky130_fd_sc_hd__o221a_1 _5402_ (.A1(_1133_),
    .A2(net535),
    .B1(_1136_),
    .B2(_1137_),
    .C1(net546),
    .X(_1140_));
 sky130_fd_sc_hd__o21ba_1 _5403_ (.A1(_1136_),
    .A2(_1139_),
    .B1_N(net547),
    .X(_0047_));
 sky130_fd_sc_hd__nor2_1 _5404_ (.A(net39),
    .B(\nco_inst.phase_accum[3] ),
    .Y(_1141_));
 sky130_fd_sc_hd__and2_1 _5405_ (.A(net39),
    .B(\nco_inst.phase_accum[3] ),
    .X(_1142_));
 sky130_fd_sc_hd__nor2_1 _5406_ (.A(_1141_),
    .B(net571),
    .Y(_1143_));
 sky130_fd_sc_hd__nand2_1 _5407_ (.A(net36),
    .B(\nco_inst.phase_accum[2] ),
    .Y(_1144_));
 sky130_fd_sc_hd__o31ai_2 _5408_ (.A1(_1133_),
    .A2(_1136_),
    .A3(_1138_),
    .B1(net538),
    .Y(_1145_));
 sky130_fd_sc_hd__xor2_1 _5409_ (.A(_1143_),
    .B(net539),
    .X(_0050_));
 sky130_fd_sc_hd__nor2_1 _5410_ (.A(net40),
    .B(\nco_inst.phase_accum[4] ),
    .Y(_1146_));
 sky130_fd_sc_hd__and2_1 _5411_ (.A(net40),
    .B(\nco_inst.phase_accum[4] ),
    .X(_1148_));
 sky130_fd_sc_hd__nor2_1 _5412_ (.A(_1146_),
    .B(net560),
    .Y(_1149_));
 sky130_fd_sc_hd__a21o_1 _5413_ (.A1(net539),
    .A2(_1143_),
    .B1(net571),
    .X(_1150_));
 sky130_fd_sc_hd__xor2_1 _5414_ (.A(_1149_),
    .B(net572),
    .X(_0051_));
 sky130_fd_sc_hd__and2_1 _5415_ (.A(net41),
    .B(\nco_inst.phase_accum[5] ),
    .X(_1151_));
 sky130_fd_sc_hd__nor2_1 _5416_ (.A(net41),
    .B(\nco_inst.phase_accum[5] ),
    .Y(_1152_));
 sky130_fd_sc_hd__or2_1 _5417_ (.A(_1151_),
    .B(net556),
    .X(_1153_));
 sky130_fd_sc_hd__a21oi_1 _5418_ (.A1(_1150_),
    .A2(_1149_),
    .B1(net560),
    .Y(_1154_));
 sky130_fd_sc_hd__xor2_1 _5419_ (.A(_1153_),
    .B(net561),
    .X(_0052_));
 sky130_fd_sc_hd__and2_1 _5420_ (.A(net42),
    .B(\nco_inst.phase_accum[6] ),
    .X(_1155_));
 sky130_fd_sc_hd__nor2_1 _5421_ (.A(net42),
    .B(\nco_inst.phase_accum[6] ),
    .Y(_1157_));
 sky130_fd_sc_hd__or2_1 _5422_ (.A(_1155_),
    .B(_1157_),
    .X(_1158_));
 sky130_fd_sc_hd__inv_2 _5423_ (.A(_1158_),
    .Y(_1159_));
 sky130_fd_sc_hd__o21bai_2 _5424_ (.A1(net556),
    .A2(_1154_),
    .B1_N(_1151_),
    .Y(_1160_));
 sky130_fd_sc_hd__xor2_1 _5425_ (.A(_1159_),
    .B(net557),
    .X(_0053_));
 sky130_fd_sc_hd__nor2_1 _5426_ (.A(net43),
    .B(\nco_inst.phase_accum[7] ),
    .Y(_1161_));
 sky130_fd_sc_hd__and2_1 _5427_ (.A(net43),
    .B(\nco_inst.phase_accum[7] ),
    .X(_1162_));
 sky130_fd_sc_hd__or2_1 _5428_ (.A(_1161_),
    .B(net674),
    .X(_1163_));
 sky130_fd_sc_hd__a21oi_2 _5429_ (.A1(net557),
    .A2(_1159_),
    .B1(_1155_),
    .Y(_1164_));
 sky130_fd_sc_hd__xor2_1 _5430_ (.A(net675),
    .B(_1164_),
    .X(_0054_));
 sky130_fd_sc_hd__xnor2_2 _5431_ (.A(net44),
    .B(\nco_inst.phase_accum[8] ),
    .Y(_1166_));
 sky130_fd_sc_hd__o21bai_2 _5432_ (.A1(_1161_),
    .A2(_1164_),
    .B1_N(net674),
    .Y(_1167_));
 sky130_fd_sc_hd__xnor2_1 _5433_ (.A(net564),
    .B(_1167_),
    .Y(_0055_));
 sky130_fd_sc_hd__nor2_1 _5434_ (.A(net45),
    .B(\nco_inst.phase_accum[9] ),
    .Y(_1168_));
 sky130_fd_sc_hd__nand2_1 _5435_ (.A(net45),
    .B(\nco_inst.phase_accum[9] ),
    .Y(_1169_));
 sky130_fd_sc_hd__and2b_1 _5436_ (.A_N(_1168_),
    .B(net634),
    .X(_1170_));
 sky130_fd_sc_hd__o21ba_1 _5437_ (.A1(_1161_),
    .A2(_1164_),
    .B1_N(_1162_),
    .X(_1171_));
 sky130_fd_sc_hd__nand2_1 _5438_ (.A(net44),
    .B(\nco_inst.phase_accum[8] ),
    .Y(_1172_));
 sky130_fd_sc_hd__o21ai_1 _5439_ (.A1(net564),
    .A2(_1171_),
    .B1(_1172_),
    .Y(_1173_));
 sky130_fd_sc_hd__xor2_1 _5440_ (.A(net635),
    .B(_1173_),
    .X(_0056_));
 sky130_fd_sc_hd__nor2_1 _5441_ (.A(net15),
    .B(\nco_inst.phase_accum[10] ),
    .Y(_1175_));
 sky130_fd_sc_hd__and2_1 _5442_ (.A(net15),
    .B(\nco_inst.phase_accum[10] ),
    .X(_1176_));
 sky130_fd_sc_hd__nor2_1 _5443_ (.A(_1175_),
    .B(net724),
    .Y(_1177_));
 sky130_fd_sc_hd__or2_1 _5444_ (.A(_1172_),
    .B(_1168_),
    .X(_1178_));
 sky130_fd_sc_hd__o311a_1 _5445_ (.A1(_1168_),
    .A2(net564),
    .A3(_1171_),
    .B1(net634),
    .C1(_1178_),
    .X(_1179_));
 sky130_fd_sc_hd__xnor2_1 _5446_ (.A(net725),
    .B(_1179_),
    .Y(_0026_));
 sky130_fd_sc_hd__xor2_1 _5447_ (.A(net16),
    .B(\nco_inst.phase_accum[11] ),
    .X(_1180_));
 sky130_fd_sc_hd__o21ba_1 _5448_ (.A1(_1175_),
    .A2(_1179_),
    .B1_N(_1176_),
    .X(_1181_));
 sky130_fd_sc_hd__xnor2_1 _5449_ (.A(net578),
    .B(_1181_),
    .Y(_0027_));
 sky130_fd_sc_hd__and4b_1 _5450_ (.A_N(_1166_),
    .B(_1170_),
    .C(_1177_),
    .D(_1180_),
    .X(_1182_));
 sky130_fd_sc_hd__o21ai_1 _5451_ (.A1(_1172_),
    .A2(_1168_),
    .B1(net634),
    .Y(_1184_));
 sky130_fd_sc_hd__a22o_1 _5452_ (.A1(net15),
    .A2(\nco_inst.phase_accum[10] ),
    .B1(net16),
    .B2(\nco_inst.phase_accum[11] ),
    .X(_1185_));
 sky130_fd_sc_hd__o21a_1 _5453_ (.A1(net16),
    .A2(\nco_inst.phase_accum[11] ),
    .B1(_1185_),
    .X(_1186_));
 sky130_fd_sc_hd__a31o_1 _5454_ (.A1(_1177_),
    .A2(_1184_),
    .A3(_1180_),
    .B1(_1186_),
    .X(_1187_));
 sky130_fd_sc_hd__a21oi_4 _5455_ (.A1(_1167_),
    .A2(_1182_),
    .B1(_1187_),
    .Y(_1188_));
 sky130_fd_sc_hd__and2_1 _5456_ (.A(net17),
    .B(\nco_inst.phase_accum[12] ),
    .X(_1189_));
 sky130_fd_sc_hd__nor2_1 _5457_ (.A(net17),
    .B(\nco_inst.phase_accum[12] ),
    .Y(_1190_));
 sky130_fd_sc_hd__nor2_1 _5458_ (.A(_1189_),
    .B(net728),
    .Y(_1191_));
 sky130_fd_sc_hd__xnor2_1 _5459_ (.A(_1188_),
    .B(net729),
    .Y(_0028_));
 sky130_fd_sc_hd__xor2_1 _5460_ (.A(net18),
    .B(\nco_inst.phase_accum[13] ),
    .X(_1192_));
 sky130_fd_sc_hd__o21ba_1 _5461_ (.A1(_1188_),
    .A2(_1190_),
    .B1_N(_1189_),
    .X(_1194_));
 sky130_fd_sc_hd__xnor2_1 _5462_ (.A(net696),
    .B(_1194_),
    .Y(_0029_));
 sky130_fd_sc_hd__or4b_1 _5463_ (.A(_1188_),
    .B(_1189_),
    .C(net728),
    .D_N(net696),
    .X(_1195_));
 sky130_fd_sc_hd__xor2_2 _5464_ (.A(net19),
    .B(net735),
    .X(_1196_));
 sky130_fd_sc_hd__a22o_1 _5465_ (.A1(net17),
    .A2(\nco_inst.phase_accum[12] ),
    .B1(net18),
    .B2(\nco_inst.phase_accum[13] ),
    .X(_1197_));
 sky130_fd_sc_hd__o21a_1 _5466_ (.A1(net18),
    .A2(\nco_inst.phase_accum[13] ),
    .B1(_1197_),
    .X(_1198_));
 sky130_fd_sc_hd__nor2_1 _5467_ (.A(_1196_),
    .B(_1198_),
    .Y(_1199_));
 sky130_fd_sc_hd__o21ai_1 _5468_ (.A1(net18),
    .A2(\nco_inst.phase_accum[13] ),
    .B1(_1197_),
    .Y(_1200_));
 sky130_fd_sc_hd__a21boi_1 _5469_ (.A1(_1195_),
    .A2(_1200_),
    .B1_N(_1196_),
    .Y(_1201_));
 sky130_fd_sc_hd__a21oi_1 _5470_ (.A1(_1195_),
    .A2(net736),
    .B1(_1201_),
    .Y(_0030_));
 sky130_fd_sc_hd__nor2_1 _5471_ (.A(net20),
    .B(\nco_inst.phase_accum[15] ),
    .Y(_1203_));
 sky130_fd_sc_hd__and2_1 _5472_ (.A(net20),
    .B(\nco_inst.phase_accum[15] ),
    .X(_1204_));
 sky130_fd_sc_hd__nor2_1 _5473_ (.A(_1203_),
    .B(_1204_),
    .Y(_1205_));
 sky130_fd_sc_hd__a21o_1 _5474_ (.A1(net19),
    .A2(\nco_inst.phase_accum[14] ),
    .B1(_1201_),
    .X(_1206_));
 sky130_fd_sc_hd__xor2_1 _5475_ (.A(_1205_),
    .B(net594),
    .X(_0031_));
 sky130_fd_sc_hd__nor2_1 _5476_ (.A(net21),
    .B(\nco_inst.phase_accum[16] ),
    .Y(_1207_));
 sky130_fd_sc_hd__nand2_1 _5477_ (.A(net21),
    .B(\nco_inst.phase_accum[16] ),
    .Y(_1208_));
 sky130_fd_sc_hd__and2b_1 _5478_ (.A_N(_1207_),
    .B(net567),
    .X(_1209_));
 sky130_fd_sc_hd__nand4_1 _5479_ (.A(_1191_),
    .B(net696),
    .C(_1196_),
    .D(_1205_),
    .Y(_1210_));
 sky130_fd_sc_hd__o211a_1 _5480_ (.A1(net20),
    .A2(\nco_inst.phase_accum[15] ),
    .B1(net19),
    .C1(\nco_inst.phase_accum[14] ),
    .X(_1211_));
 sky130_fd_sc_hd__a311o_1 _5481_ (.A1(_1196_),
    .A2(_1198_),
    .A3(_1205_),
    .B1(net706),
    .C1(_1204_),
    .X(_1213_));
 sky130_fd_sc_hd__o21bai_2 _5482_ (.A1(_1210_),
    .A2(_1188_),
    .B1_N(net707),
    .Y(_1214_));
 sky130_fd_sc_hd__xor2_1 _5483_ (.A(_1209_),
    .B(net708),
    .X(_0032_));
 sky130_fd_sc_hd__xor2_1 _5484_ (.A(net22),
    .B(\nco_inst.phase_accum[17] ),
    .X(_1215_));
 sky130_fd_sc_hd__o21ba_1 _5485_ (.A1(_1210_),
    .A2(_1188_),
    .B1_N(_1213_),
    .X(_1216_));
 sky130_fd_sc_hd__o21ai_1 _5486_ (.A1(_1207_),
    .A2(_1216_),
    .B1(net567),
    .Y(_1217_));
 sky130_fd_sc_hd__xor2_1 _5487_ (.A(_1215_),
    .B(net568),
    .X(_0033_));
 sky130_fd_sc_hd__or4bb_1 _5488_ (.A(_1207_),
    .B(_1216_),
    .C_N(_1215_),
    .D_N(_1208_),
    .X(_1218_));
 sky130_fd_sc_hd__o211a_1 _5489_ (.A1(net22),
    .A2(\nco_inst.phase_accum[17] ),
    .B1(net21),
    .C1(\nco_inst.phase_accum[16] ),
    .X(_1219_));
 sky130_fd_sc_hd__a21oi_1 _5490_ (.A1(net22),
    .A2(\nco_inst.phase_accum[17] ),
    .B1(_1219_),
    .Y(_1220_));
 sky130_fd_sc_hd__nor2_1 _5491_ (.A(net23),
    .B(\nco_inst.phase_accum[18] ),
    .Y(_1222_));
 sky130_fd_sc_hd__and2_1 _5492_ (.A(net23),
    .B(\nco_inst.phase_accum[18] ),
    .X(_1223_));
 sky130_fd_sc_hd__a211oi_1 _5493_ (.A1(_1218_),
    .A2(_1220_),
    .B1(_1222_),
    .C1(_1223_),
    .Y(_1224_));
 sky130_fd_sc_hd__o211ai_1 _5494_ (.A1(_1222_),
    .A2(_1223_),
    .B1(_1218_),
    .C1(net776),
    .Y(_1225_));
 sky130_fd_sc_hd__and2b_1 _5495_ (.A_N(_1224_),
    .B(net777),
    .X(_1226_));
 sky130_fd_sc_hd__clkbuf_1 _5496_ (.A(net778),
    .X(_0034_));
 sky130_fd_sc_hd__nor2_1 _5497_ (.A(net24),
    .B(\nco_inst.phase_accum[19] ),
    .Y(_1227_));
 sky130_fd_sc_hd__and2_1 _5498_ (.A(net24),
    .B(\nco_inst.phase_accum[19] ),
    .X(_1228_));
 sky130_fd_sc_hd__or4_1 _5499_ (.A(_1223_),
    .B(_1224_),
    .C(net688),
    .D(_1228_),
    .X(_1229_));
 sky130_fd_sc_hd__o22ai_1 _5500_ (.A1(_1223_),
    .A2(_1224_),
    .B1(net688),
    .B2(_1228_),
    .Y(_1230_));
 sky130_fd_sc_hd__nand2_1 _5501_ (.A(_1229_),
    .B(net689),
    .Y(_0035_));
 sky130_fd_sc_hd__xor2_2 _5502_ (.A(net26),
    .B(\nco_inst.phase_accum[20] ),
    .X(_1232_));
 sky130_fd_sc_hd__nor4_1 _5503_ (.A(_1222_),
    .B(_1223_),
    .C(_1227_),
    .D(_1228_),
    .Y(_1233_));
 sky130_fd_sc_hd__and3_1 _5504_ (.A(_1209_),
    .B(_1215_),
    .C(_1233_),
    .X(_1234_));
 sky130_fd_sc_hd__a21o_1 _5505_ (.A1(net22),
    .A2(\nco_inst.phase_accum[17] ),
    .B1(_1219_),
    .X(_1235_));
 sky130_fd_sc_hd__o211a_1 _5506_ (.A1(net24),
    .A2(\nco_inst.phase_accum[19] ),
    .B1(net23),
    .C1(\nco_inst.phase_accum[18] ),
    .X(_1236_));
 sky130_fd_sc_hd__a221o_1 _5507_ (.A1(net24),
    .A2(\nco_inst.phase_accum[19] ),
    .B1(_1235_),
    .B2(_1233_),
    .C1(_1236_),
    .X(_1237_));
 sky130_fd_sc_hd__a21oi_2 _5508_ (.A1(_1214_),
    .A2(_1234_),
    .B1(_1237_),
    .Y(_1238_));
 sky130_fd_sc_hd__xnor2_1 _5509_ (.A(net680),
    .B(_1238_),
    .Y(_0037_));
 sky130_fd_sc_hd__xor2_1 _5510_ (.A(net27),
    .B(\nco_inst.phase_accum[21] ),
    .X(_1239_));
 sky130_fd_sc_hd__a21o_1 _5511_ (.A1(_1214_),
    .A2(_1234_),
    .B1(_1237_),
    .X(_1241_));
 sky130_fd_sc_hd__a22oi_1 _5512_ (.A1(net26),
    .A2(\nco_inst.phase_accum[20] ),
    .B1(_1232_),
    .B2(_1241_),
    .Y(_1242_));
 sky130_fd_sc_hd__xnor2_1 _5513_ (.A(net553),
    .B(_1242_),
    .Y(_0038_));
 sky130_fd_sc_hd__and3_1 _5514_ (.A(net680),
    .B(_1241_),
    .C(net553),
    .X(_1243_));
 sky130_fd_sc_hd__xor2_1 _5515_ (.A(net28),
    .B(\nco_inst.phase_accum[22] ),
    .X(_1244_));
 sky130_fd_sc_hd__a22o_1 _5516_ (.A1(net26),
    .A2(\nco_inst.phase_accum[20] ),
    .B1(net27),
    .B2(net743),
    .X(_1245_));
 sky130_fd_sc_hd__o21a_1 _5517_ (.A1(net27),
    .A2(net743),
    .B1(_1245_),
    .X(_1246_));
 sky130_fd_sc_hd__or2_1 _5518_ (.A(_1244_),
    .B(net744),
    .X(_1247_));
 sky130_fd_sc_hd__o21a_1 _5519_ (.A1(_1243_),
    .A2(_1246_),
    .B1(_1244_),
    .X(_1248_));
 sky130_fd_sc_hd__o21ba_1 _5520_ (.A1(_1243_),
    .A2(net745),
    .B1_N(_1248_),
    .X(_0039_));
 sky130_fd_sc_hd__nor2_1 _5521_ (.A(net29),
    .B(\nco_inst.phase_accum[23] ),
    .Y(_1250_));
 sky130_fd_sc_hd__and2_1 _5522_ (.A(net29),
    .B(\nco_inst.phase_accum[23] ),
    .X(_1251_));
 sky130_fd_sc_hd__nor2_1 _5523_ (.A(_1250_),
    .B(_1251_),
    .Y(_1252_));
 sky130_fd_sc_hd__a21o_1 _5524_ (.A1(net28),
    .A2(\nco_inst.phase_accum[22] ),
    .B1(_1248_),
    .X(_1253_));
 sky130_fd_sc_hd__xor2_1 _5525_ (.A(_1252_),
    .B(net542),
    .X(_0040_));
 sky130_fd_sc_hd__nor2_1 _5526_ (.A(net460),
    .B(net30),
    .Y(_1254_));
 sky130_fd_sc_hd__nand2_1 _5527_ (.A(net460),
    .B(net30),
    .Y(_1255_));
 sky130_fd_sc_hd__and2b_1 _5528_ (.A_N(_1254_),
    .B(_1255_),
    .X(_1256_));
 sky130_fd_sc_hd__nand4_1 _5529_ (.A(net680),
    .B(net553),
    .C(_1244_),
    .D(_1252_),
    .Y(_1257_));
 sky130_fd_sc_hd__o211a_1 _5530_ (.A1(net29),
    .A2(\nco_inst.phase_accum[23] ),
    .B1(net28),
    .C1(\nco_inst.phase_accum[22] ),
    .X(_1258_));
 sky130_fd_sc_hd__a311oi_1 _5531_ (.A1(_1244_),
    .A2(_1246_),
    .A3(_1252_),
    .B1(_1258_),
    .C1(_1251_),
    .Y(_1260_));
 sky130_fd_sc_hd__o21ai_1 _5532_ (.A1(_1238_),
    .A2(_1257_),
    .B1(_1260_),
    .Y(_1261_));
 sky130_fd_sc_hd__xor2_1 _5533_ (.A(_1256_),
    .B(_1261_),
    .X(_0041_));
 sky130_fd_sc_hd__xor2_1 _5534_ (.A(net453),
    .B(net31),
    .X(_1262_));
 sky130_fd_sc_hd__o21a_1 _5535_ (.A1(_1238_),
    .A2(_1257_),
    .B1(_1260_),
    .X(_1263_));
 sky130_fd_sc_hd__o21a_1 _5536_ (.A1(_1254_),
    .A2(_1263_),
    .B1(_1255_),
    .X(_1264_));
 sky130_fd_sc_hd__xnor2_1 _5537_ (.A(_1262_),
    .B(_1264_),
    .Y(_0042_));
 sky130_fd_sc_hd__nor2_1 _5538_ (.A(net446),
    .B(net32),
    .Y(_1265_));
 sky130_fd_sc_hd__and2_1 _5539_ (.A(net447),
    .B(net32),
    .X(_1266_));
 sky130_fd_sc_hd__and3b_1 _5540_ (.A_N(_1254_),
    .B(_1262_),
    .C(_1255_),
    .X(_1267_));
 sky130_fd_sc_hd__o21a_1 _5541_ (.A1(net453),
    .A2(net31),
    .B1(net30),
    .X(_1269_));
 sky130_fd_sc_hd__a22o_1 _5542_ (.A1(net453),
    .A2(net31),
    .B1(_1269_),
    .B2(net460),
    .X(_1270_));
 sky130_fd_sc_hd__a21oi_1 _5543_ (.A1(_1261_),
    .A2(_1267_),
    .B1(_1270_),
    .Y(_1271_));
 sky130_fd_sc_hd__o21ai_1 _5544_ (.A1(_1265_),
    .A2(_1266_),
    .B1(_1271_),
    .Y(_1272_));
 sky130_fd_sc_hd__or3_1 _5545_ (.A(_1265_),
    .B(_1266_),
    .C(_1271_),
    .X(_1273_));
 sky130_fd_sc_hd__and2_1 _5546_ (.A(net803),
    .B(_1273_),
    .X(_1274_));
 sky130_fd_sc_hd__clkbuf_1 _5547_ (.A(_1274_),
    .X(_0043_));
 sky130_fd_sc_hd__xor2_1 _5548_ (.A(net435),
    .B(net33),
    .X(_1275_));
 sky130_fd_sc_hd__o21ba_1 _5549_ (.A1(_1265_),
    .A2(_1271_),
    .B1_N(_1266_),
    .X(_1276_));
 sky130_fd_sc_hd__xnor2_1 _5550_ (.A(_1275_),
    .B(_1276_),
    .Y(_0044_));
 sky130_fd_sc_hd__nand2_1 _5551_ (.A(net421),
    .B(net34),
    .Y(_1278_));
 sky130_fd_sc_hd__or2_1 _5552_ (.A(net421),
    .B(net34),
    .X(_1279_));
 sky130_fd_sc_hd__or3b_1 _5553_ (.A(_1265_),
    .B(_1266_),
    .C_N(_1275_),
    .X(_1280_));
 sky130_fd_sc_hd__o211a_1 _5554_ (.A1(net435),
    .A2(net33),
    .B1(net32),
    .C1(net447),
    .X(_1281_));
 sky130_fd_sc_hd__a21oi_1 _5555_ (.A1(net435),
    .A2(net33),
    .B1(_1281_),
    .Y(_1282_));
 sky130_fd_sc_hd__o21ai_1 _5556_ (.A1(_1280_),
    .A2(_1271_),
    .B1(_1282_),
    .Y(_1283_));
 sky130_fd_sc_hd__a21oi_1 _5557_ (.A1(_1278_),
    .A2(_1279_),
    .B1(_1283_),
    .Y(_1284_));
 sky130_fd_sc_hd__and3_1 _5558_ (.A(_1283_),
    .B(_1278_),
    .C(_1279_),
    .X(_1285_));
 sky130_fd_sc_hd__nor2_1 _5559_ (.A(net550),
    .B(_1285_),
    .Y(_0045_));
 sky130_fd_sc_hd__nor2_1 _5560_ (.A(net413),
    .B(net35),
    .Y(_1286_));
 sky130_fd_sc_hd__nand2_1 _5561_ (.A(net413),
    .B(net35),
    .Y(_1288_));
 sky130_fd_sc_hd__or2b_1 _5562_ (.A(_1286_),
    .B_N(_1288_),
    .X(_1289_));
 sky130_fd_sc_hd__a21boi_2 _5563_ (.A1(_1283_),
    .A2(_1279_),
    .B1_N(_1278_),
    .Y(_1290_));
 sky130_fd_sc_hd__xor2_1 _5564_ (.A(_1289_),
    .B(_1290_),
    .X(_0046_));
 sky130_fd_sc_hd__xor2_1 _5565_ (.A(net406),
    .B(net37),
    .X(_1291_));
 sky130_fd_sc_hd__o21ai_1 _5566_ (.A1(_1286_),
    .A2(_1290_),
    .B1(_1288_),
    .Y(_1292_));
 sky130_fd_sc_hd__xor2_1 _5567_ (.A(net714),
    .B(_1292_),
    .X(_0048_));
 sky130_fd_sc_hd__nand2_1 _5568_ (.A(net406),
    .B(net37),
    .Y(_1293_));
 sky130_fd_sc_hd__nand2_1 _5569_ (.A(_1290_),
    .B(_1288_),
    .Y(_1294_));
 sky130_fd_sc_hd__o211ai_1 _5570_ (.A1(net413),
    .A2(net35),
    .B1(_1291_),
    .C1(_1294_),
    .Y(_1295_));
 sky130_fd_sc_hd__xor2_1 _5571_ (.A(net401),
    .B(net38),
    .X(_1297_));
 sky130_fd_sc_hd__a21o_1 _5572_ (.A1(_1293_),
    .A2(_1295_),
    .B1(_1297_),
    .X(_1298_));
 sky130_fd_sc_hd__nand3_1 _5573_ (.A(_1293_),
    .B(_1295_),
    .C(_1297_),
    .Y(_1299_));
 sky130_fd_sc_hd__nand2_1 _5574_ (.A(_1298_),
    .B(net795),
    .Y(_0049_));
 sky130_fd_sc_hd__and3_1 _5575_ (.A(net237),
    .B(net380),
    .C(_0062_),
    .X(_1300_));
 sky130_fd_sc_hd__buf_2 _5576_ (.A(_1129_),
    .X(_1301_));
 sky130_fd_sc_hd__o2bb2a_1 _5577_ (.A1_N(net390),
    .A2_N(net240),
    .B1(_2982_),
    .B2(_1301_),
    .X(_1302_));
 sky130_fd_sc_hd__nor2_1 _5578_ (.A(_1300_),
    .B(_1302_),
    .Y(_0063_));
 sky130_fd_sc_hd__a22oi_2 _5579_ (.A1(net237),
    .A2(net379),
    .B1(net231),
    .B2(net391),
    .Y(_1303_));
 sky130_fd_sc_hd__nand2_1 _5580_ (.A(net245),
    .B(net367),
    .Y(_1304_));
 sky130_fd_sc_hd__a41o_1 _5581_ (.A1(net390),
    .A2(net237),
    .A3(net379),
    .A4(net231),
    .B1(_1304_),
    .X(_1306_));
 sky130_fd_sc_hd__nand4_1 _5582_ (.A(net390),
    .B(net237),
    .C(net379),
    .D(net231),
    .Y(_1307_));
 sky130_fd_sc_hd__a22o_1 _5583_ (.A1(net237),
    .A2(net379),
    .B1(net231),
    .B2(net390),
    .X(_1308_));
 sky130_fd_sc_hd__a22o_1 _5584_ (.A1(net245),
    .A2(net367),
    .B1(_1307_),
    .B2(_1308_),
    .X(_1309_));
 sky130_fd_sc_hd__o21ai_1 _5585_ (.A1(_1303_),
    .A2(_1306_),
    .B1(_1309_),
    .Y(_1310_));
 sky130_fd_sc_hd__xnor2_1 _5586_ (.A(_1300_),
    .B(_1310_),
    .Y(_0064_));
 sky130_fd_sc_hd__o211a_1 _5587_ (.A1(_1303_),
    .A2(_1306_),
    .B1(_1300_),
    .C1(_1309_),
    .X(_1311_));
 sky130_fd_sc_hd__nand4_1 _5588_ (.A(net237),
    .B(net379),
    .C(net231),
    .D(net367),
    .Y(_1312_));
 sky130_fd_sc_hd__nand2_1 _5589_ (.A(net379),
    .B(net231),
    .Y(_1313_));
 sky130_fd_sc_hd__nand2_1 _5590_ (.A(net237),
    .B(net367),
    .Y(_1314_));
 sky130_fd_sc_hd__nand2_1 _5591_ (.A(_1313_),
    .B(_1314_),
    .Y(_1316_));
 sky130_fd_sc_hd__a22o_1 _5592_ (.A1(net245),
    .A2(net356),
    .B1(_1312_),
    .B2(_1316_),
    .X(_1317_));
 sky130_fd_sc_hd__nand2_1 _5593_ (.A(net245),
    .B(net355),
    .Y(_1318_));
 sky130_fd_sc_hd__a41oi_2 _5594_ (.A1(net238),
    .A2(net379),
    .A3(net231),
    .A4(net367),
    .B1(_1318_),
    .Y(_1319_));
 sky130_fd_sc_hd__nand2_1 _5595_ (.A(_1319_),
    .B(_1316_),
    .Y(_1320_));
 sky130_fd_sc_hd__a21o_1 _5596_ (.A1(_1304_),
    .A2(_1307_),
    .B1(_1303_),
    .X(_1321_));
 sky130_fd_sc_hd__a21boi_1 _5597_ (.A1(_1317_),
    .A2(_1320_),
    .B1_N(_1321_),
    .Y(_1322_));
 sky130_fd_sc_hd__a22oi_1 _5598_ (.A1(net245),
    .A2(net356),
    .B1(_1312_),
    .B2(_1316_),
    .Y(_1323_));
 sky130_fd_sc_hd__a211oi_1 _5599_ (.A1(_1319_),
    .A2(_1316_),
    .B1(_1323_),
    .C1(_1321_),
    .Y(_1324_));
 sky130_fd_sc_hd__nor2_1 _5600_ (.A(_1322_),
    .B(_1324_),
    .Y(_1325_));
 sky130_fd_sc_hd__nand2_1 _5601_ (.A(_1311_),
    .B(_1325_),
    .Y(_1327_));
 sky130_fd_sc_hd__or2_1 _5602_ (.A(_1311_),
    .B(_1325_),
    .X(_1328_));
 sky130_fd_sc_hd__buf_4 _5603_ (.A(_3125_),
    .X(_1329_));
 sky130_fd_sc_hd__inv_2 _5604_ (.A(net227),
    .Y(_1330_));
 sky130_fd_sc_hd__buf_6 _5605_ (.A(_1330_),
    .X(_1331_));
 sky130_fd_sc_hd__buf_6 _5606_ (.A(_1331_),
    .X(_1332_));
 sky130_fd_sc_hd__o2bb2a_1 _5607_ (.A1_N(_1327_),
    .A2_N(_1328_),
    .B1(_1329_),
    .B2(_1332_),
    .X(_1333_));
 sky130_fd_sc_hd__nor2_2 _5608_ (.A(_1329_),
    .B(_1332_),
    .Y(_1334_));
 sky130_fd_sc_hd__and3_1 _5609_ (.A(_1327_),
    .B(_1328_),
    .C(_1334_),
    .X(_1335_));
 sky130_fd_sc_hd__nor2_1 _5610_ (.A(_1333_),
    .B(_1335_),
    .Y(_0065_));
 sky130_fd_sc_hd__o21ai_1 _5611_ (.A1(_1311_),
    .A2(_1325_),
    .B1(_1334_),
    .Y(_1337_));
 sky130_fd_sc_hd__nand4_2 _5612_ (.A(net238),
    .B(net233),
    .C(net367),
    .D(net355),
    .Y(_1338_));
 sky130_fd_sc_hd__nand2_1 _5613_ (.A(net232),
    .B(net368),
    .Y(_1339_));
 sky130_fd_sc_hd__nand2_1 _5614_ (.A(net240),
    .B(net355),
    .Y(_1340_));
 sky130_fd_sc_hd__nand2_1 _5615_ (.A(_1339_),
    .B(_1340_),
    .Y(_1341_));
 sky130_fd_sc_hd__a22o_1 _5616_ (.A1(net246),
    .A2(net343),
    .B1(_1338_),
    .B2(_1341_),
    .X(_1342_));
 sky130_fd_sc_hd__nand4_1 _5617_ (.A(_1341_),
    .B(net343),
    .C(net246),
    .D(_1338_),
    .Y(_1343_));
 sky130_fd_sc_hd__a22oi_1 _5618_ (.A1(net379),
    .A2(net231),
    .B1(net367),
    .B2(net237),
    .Y(_1344_));
 sky130_fd_sc_hd__o21ai_1 _5619_ (.A1(_1318_),
    .A2(_1344_),
    .B1(_1312_),
    .Y(_1345_));
 sky130_fd_sc_hd__nand3_2 _5620_ (.A(_1342_),
    .B(_1343_),
    .C(_1345_),
    .Y(_1346_));
 sky130_fd_sc_hd__nand2_1 _5621_ (.A(net245),
    .B(net343),
    .Y(_1348_));
 sky130_fd_sc_hd__a21o_1 _5622_ (.A1(_1338_),
    .A2(_1341_),
    .B1(_1348_),
    .X(_1349_));
 sky130_fd_sc_hd__o211ai_1 _5623_ (.A1(_1301_),
    .A2(_0385_),
    .B1(_1338_),
    .C1(_1341_),
    .Y(_1350_));
 sky130_fd_sc_hd__nand3b_1 _5624_ (.A_N(_1345_),
    .B(_1349_),
    .C(_1350_),
    .Y(_1351_));
 sky130_fd_sc_hd__a21o_1 _5625_ (.A1(_1316_),
    .A2(_1319_),
    .B1(_1323_),
    .X(_1352_));
 sky130_fd_sc_hd__o2bb2ai_2 _5626_ (.A1_N(_1346_),
    .A2_N(_1351_),
    .B1(_1321_),
    .B2(_1352_),
    .Y(_1353_));
 sky130_fd_sc_hd__nand3_1 _5627_ (.A(_1324_),
    .B(_1346_),
    .C(_1351_),
    .Y(_1354_));
 sky130_fd_sc_hd__inv_2 _5628_ (.A(net225),
    .Y(_1355_));
 sky130_fd_sc_hd__o22a_1 _5629_ (.A1(_2982_),
    .A2(_1332_),
    .B1(_1355_),
    .B2(_1329_),
    .X(_1356_));
 sky130_fd_sc_hd__a31o_1 _5630_ (.A1(net380),
    .A2(net225),
    .A3(_1334_),
    .B1(_1356_),
    .X(_1357_));
 sky130_fd_sc_hd__a21o_1 _5631_ (.A1(_1353_),
    .A2(_1354_),
    .B1(_1357_),
    .X(_1359_));
 sky130_fd_sc_hd__nand3_1 _5632_ (.A(_1353_),
    .B(_1354_),
    .C(_1357_),
    .Y(_1360_));
 sky130_fd_sc_hd__a22o_1 _5633_ (.A1(_1327_),
    .A2(_1337_),
    .B1(_1359_),
    .B2(_1360_),
    .X(_1361_));
 sky130_fd_sc_hd__nand4_1 _5634_ (.A(_1327_),
    .B(_1337_),
    .C(_1359_),
    .D(_1360_),
    .Y(_1362_));
 sky130_fd_sc_hd__and2_1 _5635_ (.A(_1361_),
    .B(_1362_),
    .X(_1363_));
 sky130_fd_sc_hd__clkbuf_1 _5636_ (.A(_1363_),
    .X(_0066_));
 sky130_fd_sc_hd__and2_1 _5637_ (.A(net380),
    .B(net225),
    .X(_1364_));
 sky130_fd_sc_hd__a21oi_2 _5638_ (.A1(net390),
    .A2(net215),
    .B1(_1364_),
    .Y(_1365_));
 sky130_fd_sc_hd__buf_4 _5639_ (.A(_1330_),
    .X(_1366_));
 sky130_fd_sc_hd__clkinv_4 _5640_ (.A(net214),
    .Y(_1367_));
 sky130_fd_sc_hd__nand3_2 _5641_ (.A(net390),
    .B(net380),
    .C(net221),
    .Y(_1369_));
 sky130_fd_sc_hd__o22a_1 _5642_ (.A1(_2218_),
    .A2(_1366_),
    .B1(_1367_),
    .B2(_1369_),
    .X(_1370_));
 sky130_fd_sc_hd__nand4_2 _5643_ (.A(net381),
    .B(net369),
    .C(net221),
    .D(net219),
    .Y(_1371_));
 sky130_fd_sc_hd__nand2_1 _5644_ (.A(net381),
    .B(net214),
    .Y(_1372_));
 sky130_fd_sc_hd__nand2_4 _5645_ (.A(net369),
    .B(net220),
    .Y(_1373_));
 sky130_fd_sc_hd__nand2_4 _5646_ (.A(_1372_),
    .B(_1373_),
    .Y(_1374_));
 sky130_fd_sc_hd__a2bb2oi_1 _5647_ (.A1_N(_1331_),
    .A2_N(_3134_),
    .B1(_1371_),
    .B2(_1374_),
    .Y(_1375_));
 sky130_fd_sc_hd__nand2_2 _5648_ (.A(net380),
    .B(net221),
    .Y(_1376_));
 sky130_fd_sc_hd__nand2_2 _5649_ (.A(net369),
    .B(net214),
    .Y(_1377_));
 sky130_fd_sc_hd__and2_1 _5650_ (.A(net227),
    .B(net355),
    .X(_1378_));
 sky130_fd_sc_hd__o211a_1 _5651_ (.A1(_1376_),
    .A2(_1377_),
    .B1(_1378_),
    .C1(_1374_),
    .X(_1380_));
 sky130_fd_sc_hd__o22ai_4 _5652_ (.A1(_1365_),
    .A2(_1370_),
    .B1(_1375_),
    .B2(_1380_),
    .Y(_1381_));
 sky130_fd_sc_hd__nand2_1 _5653_ (.A(net390),
    .B(net215),
    .Y(_1382_));
 sky130_fd_sc_hd__nand2_2 _5654_ (.A(_1376_),
    .B(_1382_),
    .Y(_1383_));
 sky130_fd_sc_hd__and2_1 _5655_ (.A(net368),
    .B(net227),
    .X(_1384_));
 sky130_fd_sc_hd__nand4_1 _5656_ (.A(net390),
    .B(net380),
    .C(net221),
    .D(net215),
    .Y(_1385_));
 sky130_fd_sc_hd__a21bo_1 _5657_ (.A1(_1383_),
    .A2(_1384_),
    .B1_N(_1385_),
    .X(_1386_));
 sky130_fd_sc_hd__o2bb2ai_2 _5658_ (.A1_N(_1371_),
    .A2_N(_1374_),
    .B1(_1366_),
    .B2(_3134_),
    .Y(_1387_));
 sky130_fd_sc_hd__o2111ai_4 _5659_ (.A1(_1376_),
    .A2(_1377_),
    .B1(net227),
    .C1(net355),
    .D1(_1374_),
    .Y(_1388_));
 sky130_fd_sc_hd__nand3_4 _5660_ (.A(_1386_),
    .B(_1387_),
    .C(_1388_),
    .Y(_1389_));
 sky130_fd_sc_hd__nand4_2 _5661_ (.A(_1381_),
    .B(_1389_),
    .C(net391),
    .D(net209),
    .Y(_1391_));
 sky130_fd_sc_hd__inv_2 _5662_ (.A(_1391_),
    .Y(_1392_));
 sky130_fd_sc_hd__inv_6 _5663_ (.A(net208),
    .Y(_1393_));
 sky130_fd_sc_hd__clkbuf_4 _5664_ (.A(_1393_),
    .X(_1394_));
 sky130_fd_sc_hd__o2bb2a_1 _5665_ (.A1_N(_1381_),
    .A2_N(_1389_),
    .B1(_1329_),
    .B2(_1394_),
    .X(_1395_));
 sky130_fd_sc_hd__nor2_1 _5666_ (.A(_1392_),
    .B(_1395_),
    .Y(_1396_));
 sky130_fd_sc_hd__a2111o_1 _5667_ (.A1(_2218_),
    .A2(net219),
    .B1(_1376_),
    .C1(_1332_),
    .D1(_1329_),
    .X(_1397_));
 sky130_fd_sc_hd__nand2_1 _5668_ (.A(net232),
    .B(net343),
    .Y(_1398_));
 sky130_fd_sc_hd__nand2_1 _5669_ (.A(net238),
    .B(net328),
    .Y(_1399_));
 sky130_fd_sc_hd__nand2_1 _5670_ (.A(_1398_),
    .B(_1399_),
    .Y(_1400_));
 sky130_fd_sc_hd__nand4_4 _5671_ (.A(net239),
    .B(net232),
    .C(net343),
    .D(net329),
    .Y(_1402_));
 sky130_fd_sc_hd__a22o_1 _5672_ (.A1(net245),
    .A2(net316),
    .B1(_1400_),
    .B2(_1402_),
    .X(_1403_));
 sky130_fd_sc_hd__nand2_1 _5673_ (.A(net247),
    .B(net328),
    .Y(_1404_));
 sky130_fd_sc_hd__a22oi_1 _5674_ (.A1(net233),
    .A2(net355),
    .B1(net343),
    .B2(net240),
    .Y(_1405_));
 sky130_fd_sc_hd__nand4_2 _5675_ (.A(net240),
    .B(net233),
    .C(net355),
    .D(net344),
    .Y(_1406_));
 sky130_fd_sc_hd__o21ai_2 _5676_ (.A1(_1404_),
    .A2(_1405_),
    .B1(_1406_),
    .Y(_1407_));
 sky130_fd_sc_hd__nand4_2 _5677_ (.A(_1400_),
    .B(_1402_),
    .C(net245),
    .D(net316),
    .Y(_1408_));
 sky130_fd_sc_hd__nand3_2 _5678_ (.A(_1403_),
    .B(_1407_),
    .C(_1408_),
    .Y(_1409_));
 sky130_fd_sc_hd__nand2_1 _5679_ (.A(net246),
    .B(net316),
    .Y(_1410_));
 sky130_fd_sc_hd__a21o_1 _5680_ (.A1(_1400_),
    .A2(_1402_),
    .B1(_1410_),
    .X(_1411_));
 sky130_fd_sc_hd__o211ai_1 _5681_ (.A1(_1301_),
    .A2(net96),
    .B1(_1400_),
    .C1(_1402_),
    .Y(_1413_));
 sky130_fd_sc_hd__nand3b_2 _5682_ (.A_N(_1407_),
    .B(_1411_),
    .C(_1413_),
    .Y(_1414_));
 sky130_fd_sc_hd__buf_4 _5683_ (.A(_1367_),
    .X(_1415_));
 sky130_fd_sc_hd__o2111ai_4 _5684_ (.A1(_1415_),
    .A2(_1369_),
    .B1(net368),
    .C1(_1383_),
    .D1(net227),
    .Y(_1416_));
 sky130_fd_sc_hd__nand4b_4 _5685_ (.A_N(_1397_),
    .B(_1409_),
    .C(_1414_),
    .D(_1416_),
    .Y(_1417_));
 sky130_fd_sc_hd__and3_1 _5686_ (.A(_1383_),
    .B(_1384_),
    .C(_1385_),
    .X(_1418_));
 sky130_fd_sc_hd__o2bb2ai_2 _5687_ (.A1_N(_1409_),
    .A2_N(_1414_),
    .B1(_1418_),
    .B2(_1397_),
    .Y(_1419_));
 sky130_fd_sc_hd__nand2_1 _5688_ (.A(net233),
    .B(net355),
    .Y(_1420_));
 sky130_fd_sc_hd__nand2_1 _5689_ (.A(net240),
    .B(net343),
    .Y(_1421_));
 sky130_fd_sc_hd__nand2_1 _5690_ (.A(_1420_),
    .B(_1421_),
    .Y(_1422_));
 sky130_fd_sc_hd__and4_1 _5691_ (.A(_1422_),
    .B(net328),
    .C(net247),
    .D(_1406_),
    .X(_1424_));
 sky130_fd_sc_hd__a21boi_1 _5692_ (.A1(_1348_),
    .A2(_1338_),
    .B1_N(_1341_),
    .Y(_1425_));
 sky130_fd_sc_hd__o2bb2ai_1 _5693_ (.A1_N(_1406_),
    .A2_N(_1422_),
    .B1(_1129_),
    .B2(_3441_),
    .Y(_1426_));
 sky130_fd_sc_hd__nand2_1 _5694_ (.A(_1425_),
    .B(_1426_),
    .Y(_1427_));
 sky130_fd_sc_hd__o2bb2ai_1 _5695_ (.A1_N(_1417_),
    .A2_N(_1419_),
    .B1(_1424_),
    .B2(_1427_),
    .Y(_1428_));
 sky130_fd_sc_hd__o2111ai_1 _5696_ (.A1(_1340_),
    .A2(_1398_),
    .B1(net250),
    .C1(net328),
    .D1(_1422_),
    .Y(_1429_));
 sky130_fd_sc_hd__and3_1 _5697_ (.A(_1425_),
    .B(_1426_),
    .C(_1429_),
    .X(_1430_));
 sky130_fd_sc_hd__nand3_1 _5698_ (.A(_1419_),
    .B(_1430_),
    .C(_1417_),
    .Y(_1431_));
 sky130_fd_sc_hd__nand3_2 _5699_ (.A(_1396_),
    .B(_1428_),
    .C(_1431_),
    .Y(_1432_));
 sky130_fd_sc_hd__a21oi_1 _5700_ (.A1(_1426_),
    .A2(_1429_),
    .B1(_1425_),
    .Y(_1433_));
 sky130_fd_sc_hd__nor3_1 _5701_ (.A(_1346_),
    .B(_1433_),
    .C(_1430_),
    .Y(_1435_));
 sky130_fd_sc_hd__a22o_1 _5702_ (.A1(net367),
    .A2(net227),
    .B1(_1385_),
    .B2(_1383_),
    .X(_1436_));
 sky130_fd_sc_hd__a22oi_2 _5703_ (.A1(_1334_),
    .A2(_1364_),
    .B1(_1436_),
    .B2(_1416_),
    .Y(_1437_));
 sky130_fd_sc_hd__and4_1 _5704_ (.A(_1436_),
    .B(_1416_),
    .C(_1334_),
    .D(_1364_),
    .X(_1438_));
 sky130_fd_sc_hd__o21a_1 _5705_ (.A1(_1433_),
    .A2(_1430_),
    .B1(_1346_),
    .X(_1439_));
 sky130_fd_sc_hd__nor4_1 _5706_ (.A(_1435_),
    .B(_1437_),
    .C(_1438_),
    .D(_1439_),
    .Y(_1440_));
 sky130_fd_sc_hd__o211ai_1 _5707_ (.A1(_1424_),
    .A2(_1427_),
    .B1(_1417_),
    .C1(_1419_),
    .Y(_1441_));
 sky130_fd_sc_hd__a41o_1 _5708_ (.A1(net247),
    .A2(net328),
    .A3(_1406_),
    .A4(_1422_),
    .B1(_1427_),
    .X(_1442_));
 sky130_fd_sc_hd__a21o_1 _5709_ (.A1(_1417_),
    .A2(_1419_),
    .B1(_1442_),
    .X(_1443_));
 sky130_fd_sc_hd__o211ai_2 _5710_ (.A1(_1392_),
    .A2(_1395_),
    .B1(_1441_),
    .C1(_1443_),
    .Y(_1444_));
 sky130_fd_sc_hd__o21a_1 _5711_ (.A1(_1435_),
    .A2(_1440_),
    .B1(_1444_),
    .X(_1446_));
 sky130_fd_sc_hd__a211o_1 _5712_ (.A1(_1444_),
    .A2(_1432_),
    .B1(_1435_),
    .C1(_1440_),
    .X(_1447_));
 sky130_fd_sc_hd__a21bo_1 _5713_ (.A1(_1432_),
    .A2(_1446_),
    .B1_N(_1447_),
    .X(_1448_));
 sky130_fd_sc_hd__nand2_1 _5714_ (.A(_1354_),
    .B(_1357_),
    .Y(_1449_));
 sky130_fd_sc_hd__o22ai_1 _5715_ (.A1(_1437_),
    .A2(_1438_),
    .B1(_1439_),
    .B2(_1435_),
    .Y(_1450_));
 sky130_fd_sc_hd__nor2_1 _5716_ (.A(_1437_),
    .B(_1438_),
    .Y(_1451_));
 sky130_fd_sc_hd__o21ai_1 _5717_ (.A1(_1433_),
    .A2(_1430_),
    .B1(_1346_),
    .Y(_1452_));
 sky130_fd_sc_hd__nand3b_1 _5718_ (.A_N(_1435_),
    .B(_1451_),
    .C(_1452_),
    .Y(_1453_));
 sky130_fd_sc_hd__a22oi_1 _5719_ (.A1(_1353_),
    .A2(_1449_),
    .B1(_1450_),
    .B2(_1453_),
    .Y(_1454_));
 sky130_fd_sc_hd__nand4_1 _5720_ (.A(_1353_),
    .B(_1453_),
    .C(_1449_),
    .D(_1450_),
    .Y(_1455_));
 sky130_fd_sc_hd__o21ai_1 _5721_ (.A1(_1454_),
    .A2(_1361_),
    .B1(_1455_),
    .Y(_1457_));
 sky130_fd_sc_hd__xnor2_1 _5722_ (.A(_1448_),
    .B(_1457_),
    .Y(_0101_));
 sky130_fd_sc_hd__a22oi_1 _5723_ (.A1(net232),
    .A2(net343),
    .B1(net329),
    .B2(net239),
    .Y(_1458_));
 sky130_fd_sc_hd__a21oi_2 _5724_ (.A1(_1410_),
    .A2(_1402_),
    .B1(_1458_),
    .Y(_1459_));
 sky130_fd_sc_hd__nand2_1 _5725_ (.A(net232),
    .B(net328),
    .Y(_1460_));
 sky130_fd_sc_hd__nand2_1 _5726_ (.A(net240),
    .B(net316),
    .Y(_1461_));
 sky130_fd_sc_hd__nand2_1 _5727_ (.A(_1460_),
    .B(_1461_),
    .Y(_1462_));
 sky130_fd_sc_hd__nand4_2 _5728_ (.A(net239),
    .B(net232),
    .C(net328),
    .D(net316),
    .Y(_1463_));
 sky130_fd_sc_hd__a22o_1 _5729_ (.A1(net246),
    .A2(net306),
    .B1(_1462_),
    .B2(_1463_),
    .X(_1464_));
 sky130_fd_sc_hd__nand4_1 _5730_ (.A(_1462_),
    .B(_1463_),
    .C(net246),
    .D(net306),
    .Y(_1465_));
 sky130_fd_sc_hd__nand3_2 _5731_ (.A(_1459_),
    .B(_1464_),
    .C(_1465_),
    .Y(_1467_));
 sky130_fd_sc_hd__nand2_1 _5732_ (.A(net246),
    .B(net306),
    .Y(_1468_));
 sky130_fd_sc_hd__a21o_1 _5733_ (.A1(_1462_),
    .A2(_1463_),
    .B1(_1468_),
    .X(_1469_));
 sky130_fd_sc_hd__o211ai_1 _5734_ (.A1(_1301_),
    .A2(_2973_),
    .B1(_1462_),
    .C1(_1463_),
    .Y(_1470_));
 sky130_fd_sc_hd__nand3b_1 _5735_ (.A_N(_1459_),
    .B(_1469_),
    .C(_1470_),
    .Y(_1471_));
 sky130_fd_sc_hd__nand3b_2 _5736_ (.A_N(_1389_),
    .B(_1467_),
    .C(_1471_),
    .Y(_1472_));
 sky130_fd_sc_hd__inv_2 _5737_ (.A(_1472_),
    .Y(_1473_));
 sky130_fd_sc_hd__nand3b_1 _5738_ (.A_N(_1370_),
    .B(_1387_),
    .C(_1388_),
    .Y(_1474_));
 sky130_fd_sc_hd__o2bb2ai_2 _5739_ (.A1_N(_1467_),
    .A2_N(_1471_),
    .B1(_1365_),
    .B2(_1474_),
    .Y(_1475_));
 sky130_fd_sc_hd__and3_1 _5740_ (.A(_1403_),
    .B(_1407_),
    .C(_1408_),
    .X(_1476_));
 sky130_fd_sc_hd__nand2_1 _5741_ (.A(_1475_),
    .B(_1476_),
    .Y(_1478_));
 sky130_fd_sc_hd__a21o_1 _5742_ (.A1(_1475_),
    .A2(_1472_),
    .B1(_1476_),
    .X(_1479_));
 sky130_fd_sc_hd__o21ai_1 _5743_ (.A1(_1473_),
    .A2(_1478_),
    .B1(_1479_),
    .Y(_1480_));
 sky130_fd_sc_hd__nand2_1 _5744_ (.A(net356),
    .B(net220),
    .Y(_1481_));
 sky130_fd_sc_hd__nand2_2 _5745_ (.A(net356),
    .B(net214),
    .Y(_1482_));
 sky130_fd_sc_hd__o2bb2ai_1 _5746_ (.A1_N(_1377_),
    .A2_N(_1481_),
    .B1(_1482_),
    .B2(_1373_),
    .Y(_1483_));
 sky130_fd_sc_hd__o21ai_2 _5747_ (.A1(_1331_),
    .A2(_0385_),
    .B1(_1483_),
    .Y(_1484_));
 sky130_fd_sc_hd__o2bb2ai_2 _5748_ (.A1_N(_1378_),
    .A2_N(_1374_),
    .B1(_1377_),
    .B2(_1376_),
    .Y(_1485_));
 sky130_fd_sc_hd__and2_1 _5749_ (.A(net226),
    .B(net344),
    .X(_1486_));
 sky130_fd_sc_hd__a22o_1 _5750_ (.A1(net356),
    .A2(net220),
    .B1(net214),
    .B2(net369),
    .X(_1487_));
 sky130_fd_sc_hd__o211ai_4 _5751_ (.A1(_1373_),
    .A2(_1482_),
    .B1(_1486_),
    .C1(_1487_),
    .Y(_1489_));
 sky130_fd_sc_hd__nand3_4 _5752_ (.A(_1484_),
    .B(_1485_),
    .C(_1489_),
    .Y(_1490_));
 sky130_fd_sc_hd__nand2_1 _5753_ (.A(net226),
    .B(net344),
    .Y(_1491_));
 sky130_fd_sc_hd__o21ai_2 _5754_ (.A1(_1373_),
    .A2(_1482_),
    .B1(_1491_),
    .Y(_1492_));
 sky130_fd_sc_hd__a22oi_4 _5755_ (.A1(net356),
    .A2(net220),
    .B1(net214),
    .B2(net369),
    .Y(_1493_));
 sky130_fd_sc_hd__a21boi_2 _5756_ (.A1(_1374_),
    .A2(_1378_),
    .B1_N(_1371_),
    .Y(_1494_));
 sky130_fd_sc_hd__nand2_1 _5757_ (.A(_1483_),
    .B(_1486_),
    .Y(_1495_));
 sky130_fd_sc_hd__o211ai_4 _5758_ (.A1(_1492_),
    .A2(_1493_),
    .B1(_1494_),
    .C1(_1495_),
    .Y(_1496_));
 sky130_fd_sc_hd__and4_2 _5759_ (.A(net392),
    .B(net378),
    .C(net208),
    .D(net201),
    .X(_1497_));
 sky130_fd_sc_hd__nand2_1 _5760_ (.A(net391),
    .B(net202),
    .Y(_1498_));
 sky130_fd_sc_hd__o21a_1 _5761_ (.A1(_2982_),
    .A2(_1393_),
    .B1(_1498_),
    .X(_1500_));
 sky130_fd_sc_hd__o2bb2ai_2 _5762_ (.A1_N(_1490_),
    .A2_N(_1496_),
    .B1(_1497_),
    .B2(_1500_),
    .Y(_1501_));
 sky130_fd_sc_hd__nor2_2 _5763_ (.A(_3125_),
    .B(_1393_),
    .Y(_1502_));
 sky130_fd_sc_hd__and2_1 _5764_ (.A(net381),
    .B(net202),
    .X(_1503_));
 sky130_fd_sc_hd__a21oi_1 _5765_ (.A1(_1502_),
    .A2(_1503_),
    .B1(_1500_),
    .Y(_1504_));
 sky130_fd_sc_hd__nand3_2 _5766_ (.A(_1490_),
    .B(_1496_),
    .C(_1504_),
    .Y(_1505_));
 sky130_fd_sc_hd__nand2_1 _5767_ (.A(_1501_),
    .B(_1505_),
    .Y(_1506_));
 sky130_fd_sc_hd__or2_1 _5768_ (.A(_1391_),
    .B(_1506_),
    .X(_1507_));
 sky130_fd_sc_hd__a32o_1 _5769_ (.A1(_1502_),
    .A2(_1381_),
    .A3(_1389_),
    .B1(_1501_),
    .B2(_1505_),
    .X(_1508_));
 sky130_fd_sc_hd__nand3_2 _5770_ (.A(_1480_),
    .B(_1507_),
    .C(_1508_),
    .Y(_1509_));
 sky130_fd_sc_hd__a32oi_4 _5771_ (.A1(_1502_),
    .A2(_1381_),
    .A3(_1389_),
    .B1(_1501_),
    .B2(_1505_),
    .Y(_1511_));
 sky130_fd_sc_hd__nor2_1 _5772_ (.A(_1391_),
    .B(_1506_),
    .Y(_1512_));
 sky130_fd_sc_hd__o221ai_4 _5773_ (.A1(_1478_),
    .A2(_1473_),
    .B1(_1511_),
    .B2(_1512_),
    .C1(_1479_),
    .Y(_1513_));
 sky130_fd_sc_hd__a21o_1 _5774_ (.A1(_1509_),
    .A2(_1513_),
    .B1(_1432_),
    .X(_1514_));
 sky130_fd_sc_hd__nand3_1 _5775_ (.A(_1432_),
    .B(_1509_),
    .C(_1513_),
    .Y(_1515_));
 sky130_fd_sc_hd__a21bo_1 _5776_ (.A1(_1430_),
    .A2(_1419_),
    .B1_N(_1417_),
    .X(_1516_));
 sky130_fd_sc_hd__a21o_1 _5777_ (.A1(_1514_),
    .A2(_1515_),
    .B1(_1516_),
    .X(_1517_));
 sky130_fd_sc_hd__nand3_1 _5778_ (.A(_1514_),
    .B(_1515_),
    .C(_1516_),
    .Y(_1518_));
 sky130_fd_sc_hd__a22o_1 _5779_ (.A1(_1432_),
    .A2(_1446_),
    .B1(_1447_),
    .B2(_1457_),
    .X(_1519_));
 sky130_fd_sc_hd__a21oi_1 _5780_ (.A1(_1517_),
    .A2(_1518_),
    .B1(_1519_),
    .Y(_1520_));
 sky130_fd_sc_hd__nand3_1 _5781_ (.A(_1519_),
    .B(_1517_),
    .C(_1518_),
    .Y(_1522_));
 sky130_fd_sc_hd__and2b_1 _5782_ (.A_N(_1520_),
    .B(_1522_),
    .X(_1523_));
 sky130_fd_sc_hd__clkbuf_1 _5783_ (.A(_1523_),
    .X(_0102_));
 sky130_fd_sc_hd__a22oi_1 _5784_ (.A1(net232),
    .A2(net328),
    .B1(net316),
    .B2(net239),
    .Y(_1524_));
 sky130_fd_sc_hd__a21oi_2 _5785_ (.A1(_1463_),
    .A2(_1468_),
    .B1(_1524_),
    .Y(_1525_));
 sky130_fd_sc_hd__nand4_2 _5786_ (.A(net240),
    .B(net233),
    .C(net317),
    .D(net306),
    .Y(_1526_));
 sky130_fd_sc_hd__nand2_1 _5787_ (.A(net235),
    .B(net316),
    .Y(_1527_));
 sky130_fd_sc_hd__nand2_2 _5788_ (.A(net242),
    .B(net306),
    .Y(_1528_));
 sky130_fd_sc_hd__nand2_2 _5789_ (.A(_1527_),
    .B(_1528_),
    .Y(_1529_));
 sky130_fd_sc_hd__nand2_1 _5790_ (.A(net299),
    .B(net247),
    .Y(_1530_));
 sky130_fd_sc_hd__a21o_1 _5791_ (.A1(_1526_),
    .A2(_1529_),
    .B1(_1530_),
    .X(_1532_));
 sky130_fd_sc_hd__nand2_2 _5792_ (.A(net233),
    .B(net306),
    .Y(_1533_));
 sky130_fd_sc_hd__o221ai_2 _5793_ (.A1(_3022_),
    .A2(_1129_),
    .B1(_1461_),
    .B2(_1533_),
    .C1(_1529_),
    .Y(_1534_));
 sky130_fd_sc_hd__nand3b_2 _5794_ (.A_N(_1525_),
    .B(_1532_),
    .C(_1534_),
    .Y(_1535_));
 sky130_fd_sc_hd__a22o_1 _5795_ (.A1(net299),
    .A2(net247),
    .B1(_1526_),
    .B2(_1529_),
    .X(_1536_));
 sky130_fd_sc_hd__o2111ai_1 _5796_ (.A1(_1461_),
    .A2(_1533_),
    .B1(net299),
    .C1(net247),
    .D1(_1529_),
    .Y(_1537_));
 sky130_fd_sc_hd__nand3_2 _5797_ (.A(_1536_),
    .B(_1537_),
    .C(_1525_),
    .Y(_1538_));
 sky130_fd_sc_hd__nand2_1 _5798_ (.A(_1535_),
    .B(_1538_),
    .Y(_1539_));
 sky130_fd_sc_hd__nor2_2 _5799_ (.A(_1490_),
    .B(_1539_),
    .Y(_1540_));
 sky130_fd_sc_hd__a21o_1 _5800_ (.A1(_1490_),
    .A2(_1539_),
    .B1(_1467_),
    .X(_1541_));
 sky130_fd_sc_hd__nor2_1 _5801_ (.A(_1540_),
    .B(_1541_),
    .Y(_1543_));
 sky130_fd_sc_hd__and2_1 _5802_ (.A(_1464_),
    .B(_1465_),
    .X(_1544_));
 sky130_fd_sc_hd__a32oi_2 _5803_ (.A1(_1485_),
    .A2(_1489_),
    .A3(_1484_),
    .B1(_1535_),
    .B2(_1538_),
    .Y(_1545_));
 sky130_fd_sc_hd__o2bb2a_1 _5804_ (.A1_N(_1544_),
    .A2_N(_1459_),
    .B1(_1545_),
    .B2(_1540_),
    .X(_1546_));
 sky130_fd_sc_hd__and4_1 _5805_ (.A(net391),
    .B(net381),
    .C(net201),
    .D(net195),
    .X(_1547_));
 sky130_fd_sc_hd__a22oi_4 _5806_ (.A1(net381),
    .A2(net202),
    .B1(net200),
    .B2(net391),
    .Y(_1548_));
 sky130_fd_sc_hd__a211oi_2 _5807_ (.A1(net369),
    .A2(net209),
    .B1(_1547_),
    .C1(_1548_),
    .Y(_1549_));
 sky130_fd_sc_hd__o211a_1 _5808_ (.A1(_1547_),
    .A2(_1548_),
    .B1(net369),
    .C1(net209),
    .X(_1550_));
 sky130_fd_sc_hd__nand2_1 _5809_ (.A(_1502_),
    .B(_1503_),
    .Y(_1551_));
 sky130_fd_sc_hd__nand2_1 _5810_ (.A(net220),
    .B(net344),
    .Y(_1552_));
 sky130_fd_sc_hd__nand2_2 _5811_ (.A(_1482_),
    .B(_1552_),
    .Y(_1554_));
 sky130_fd_sc_hd__nand4_4 _5812_ (.A(net354),
    .B(net220),
    .C(net342),
    .D(net214),
    .Y(_1555_));
 sky130_fd_sc_hd__nand2_1 _5813_ (.A(_1554_),
    .B(_1555_),
    .Y(_1556_));
 sky130_fd_sc_hd__and2_1 _5814_ (.A(net226),
    .B(net331),
    .X(_1557_));
 sky130_fd_sc_hd__nand2_1 _5815_ (.A(_1556_),
    .B(_1557_),
    .Y(_1558_));
 sky130_fd_sc_hd__o211ai_2 _5816_ (.A1(_1331_),
    .A2(_3441_),
    .B1(_1554_),
    .C1(_1555_),
    .Y(_1559_));
 sky130_fd_sc_hd__nand3_4 _5817_ (.A(_1551_),
    .B(_1558_),
    .C(_1559_),
    .Y(_1560_));
 sky130_fd_sc_hd__a21o_1 _5818_ (.A1(_1554_),
    .A2(_1555_),
    .B1(_1557_),
    .X(_1561_));
 sky130_fd_sc_hd__nand4_2 _5819_ (.A(_1554_),
    .B(_1555_),
    .C(net226),
    .D(net331),
    .Y(_1562_));
 sky130_fd_sc_hd__nand3_4 _5820_ (.A(_1561_),
    .B(_1562_),
    .C(_1497_),
    .Y(_1563_));
 sky130_fd_sc_hd__nand4_2 _5821_ (.A(_1487_),
    .B(_1492_),
    .C(_1560_),
    .D(_1563_),
    .Y(_1565_));
 sky130_fd_sc_hd__a2bb2o_1 _5822_ (.A1_N(_1373_),
    .A2_N(_1482_),
    .B1(_1486_),
    .B2(_1487_),
    .X(_1566_));
 sky130_fd_sc_hd__a21o_1 _5823_ (.A1(_1560_),
    .A2(_1563_),
    .B1(_1566_),
    .X(_1567_));
 sky130_fd_sc_hd__o211ai_4 _5824_ (.A1(_1549_),
    .A2(_1550_),
    .B1(_1565_),
    .C1(_1567_),
    .Y(_1568_));
 sky130_fd_sc_hd__and3_1 _5825_ (.A(_1490_),
    .B(_1496_),
    .C(_1504_),
    .X(_1569_));
 sky130_fd_sc_hd__nand2_1 _5826_ (.A(_1560_),
    .B(_1563_),
    .Y(_1570_));
 sky130_fd_sc_hd__nand2_1 _5827_ (.A(_1570_),
    .B(_1566_),
    .Y(_1571_));
 sky130_fd_sc_hd__o32a_1 _5828_ (.A1(_1355_),
    .A2(_1415_),
    .A3(_0133_),
    .B1(_1491_),
    .B2(_1493_),
    .X(_1572_));
 sky130_fd_sc_hd__nand3_2 _5829_ (.A(_1560_),
    .B(_1563_),
    .C(_1572_),
    .Y(_1573_));
 sky130_fd_sc_hd__nor2_1 _5830_ (.A(_1549_),
    .B(_1550_),
    .Y(_1574_));
 sky130_fd_sc_hd__nand3_2 _5831_ (.A(_1571_),
    .B(_1573_),
    .C(_1574_),
    .Y(_1576_));
 sky130_fd_sc_hd__and3_1 _5832_ (.A(_1568_),
    .B(_1569_),
    .C(_1576_),
    .X(_1577_));
 sky130_fd_sc_hd__a21oi_1 _5833_ (.A1(_1576_),
    .A2(_1568_),
    .B1(_1569_),
    .Y(_1578_));
 sky130_fd_sc_hd__o22ai_1 _5834_ (.A1(_1543_),
    .A2(_1546_),
    .B1(_1577_),
    .B2(_1578_),
    .Y(_1579_));
 sky130_fd_sc_hd__nand3_1 _5835_ (.A(_1475_),
    .B(_1472_),
    .C(_1476_),
    .Y(_1580_));
 sky130_fd_sc_hd__a31o_1 _5836_ (.A1(_1479_),
    .A2(_1580_),
    .A3(_1508_),
    .B1(_1512_),
    .X(_1581_));
 sky130_fd_sc_hd__o2bb2ai_1 _5837_ (.A1_N(_1544_),
    .A2_N(_1459_),
    .B1(_1545_),
    .B2(_1540_),
    .Y(_1582_));
 sky130_fd_sc_hd__nand3_2 _5838_ (.A(_1568_),
    .B(_1569_),
    .C(_1576_),
    .Y(_1583_));
 sky130_fd_sc_hd__nand2_1 _5839_ (.A(_1490_),
    .B(_1496_),
    .Y(_1584_));
 sky130_fd_sc_hd__a31o_1 _5840_ (.A1(net391),
    .A2(net209),
    .A3(_1503_),
    .B1(_1500_),
    .X(_1585_));
 sky130_fd_sc_hd__o2bb2ai_2 _5841_ (.A1_N(_1576_),
    .A2_N(_1568_),
    .B1(_1584_),
    .B2(_1585_),
    .Y(_1587_));
 sky130_fd_sc_hd__o2111ai_2 _5842_ (.A1(_1540_),
    .A2(_1541_),
    .B1(_1582_),
    .C1(_1583_),
    .D1(_1587_),
    .Y(_1588_));
 sky130_fd_sc_hd__nand3_2 _5843_ (.A(_1579_),
    .B(_1581_),
    .C(_1588_),
    .Y(_1589_));
 sky130_fd_sc_hd__o21a_1 _5844_ (.A1(_1511_),
    .A2(_1480_),
    .B1(_1507_),
    .X(_1590_));
 sky130_fd_sc_hd__o21ai_1 _5845_ (.A1(_1540_),
    .A2(_1541_),
    .B1(_1582_),
    .Y(_1591_));
 sky130_fd_sc_hd__a21o_1 _5846_ (.A1(_1583_),
    .A2(_1587_),
    .B1(_1591_),
    .X(_1592_));
 sky130_fd_sc_hd__o211ai_2 _5847_ (.A1(_1543_),
    .A2(_1546_),
    .B1(_1583_),
    .C1(_1587_),
    .Y(_1593_));
 sky130_fd_sc_hd__nand3_4 _5848_ (.A(_1590_),
    .B(_1592_),
    .C(_1593_),
    .Y(_1594_));
 sky130_fd_sc_hd__nor2_1 _5849_ (.A(_1476_),
    .B(_1473_),
    .Y(_1595_));
 sky130_fd_sc_hd__inv_2 _5850_ (.A(_1475_),
    .Y(_1596_));
 sky130_fd_sc_hd__o2bb2ai_2 _5851_ (.A1_N(_1589_),
    .A2_N(_1594_),
    .B1(_1595_),
    .B2(_1596_),
    .Y(_1598_));
 sky130_fd_sc_hd__a41o_2 _5852_ (.A1(_1408_),
    .A2(_1403_),
    .A3(_1475_),
    .A4(_1407_),
    .B1(_1473_),
    .X(_1599_));
 sky130_fd_sc_hd__nand3_1 _5853_ (.A(_1589_),
    .B(_1594_),
    .C(_1599_),
    .Y(_1600_));
 sky130_fd_sc_hd__a21oi_1 _5854_ (.A1(_1509_),
    .A2(_1513_),
    .B1(_1432_),
    .Y(_1601_));
 sky130_fd_sc_hd__a21o_1 _5855_ (.A1(_1515_),
    .A2(_1516_),
    .B1(_1601_),
    .X(_1602_));
 sky130_fd_sc_hd__a21oi_1 _5856_ (.A1(_1598_),
    .A2(_1600_),
    .B1(_1602_),
    .Y(_1603_));
 sky130_fd_sc_hd__nand3_1 _5857_ (.A(_1598_),
    .B(_1600_),
    .C(_1602_),
    .Y(_1604_));
 sky130_fd_sc_hd__a21oi_1 _5858_ (.A1(_1522_),
    .A2(_1604_),
    .B1(_1603_),
    .Y(_1605_));
 sky130_fd_sc_hd__a21oi_1 _5859_ (.A1(_1522_),
    .A2(_1603_),
    .B1(_1605_),
    .Y(_0103_));
 sky130_fd_sc_hd__a21boi_4 _5860_ (.A1(_1594_),
    .A2(_1599_),
    .B1_N(_1589_),
    .Y(_1606_));
 sky130_fd_sc_hd__nand2_2 _5861_ (.A(net378),
    .B(net195),
    .Y(_1608_));
 sky130_fd_sc_hd__nand2_1 _5862_ (.A(net369),
    .B(net208),
    .Y(_1609_));
 sky130_fd_sc_hd__o21a_1 _5863_ (.A1(_1498_),
    .A2(_1608_),
    .B1(_1609_),
    .X(_1610_));
 sky130_fd_sc_hd__nand2_1 _5864_ (.A(net344),
    .B(net215),
    .Y(_1611_));
 sky130_fd_sc_hd__nand2_2 _5865_ (.A(net221),
    .B(net329),
    .Y(_1612_));
 sky130_fd_sc_hd__nand2_2 _5866_ (.A(_1611_),
    .B(_1612_),
    .Y(_1613_));
 sky130_fd_sc_hd__nand4_4 _5867_ (.A(net221),
    .B(net344),
    .C(net215),
    .D(net329),
    .Y(_1614_));
 sky130_fd_sc_hd__o211ai_2 _5868_ (.A1(_1366_),
    .A2(_1782_),
    .B1(_1613_),
    .C1(_1614_),
    .Y(_1615_));
 sky130_fd_sc_hd__nand2_1 _5869_ (.A(net228),
    .B(net317),
    .Y(_1616_));
 sky130_fd_sc_hd__a21o_1 _5870_ (.A1(_1613_),
    .A2(_1614_),
    .B1(_1616_),
    .X(_1617_));
 sky130_fd_sc_hd__o211ai_4 _5871_ (.A1(_1548_),
    .A2(_1610_),
    .B1(_1615_),
    .C1(_1617_),
    .Y(_1619_));
 sky130_fd_sc_hd__a22o_1 _5872_ (.A1(net226),
    .A2(net317),
    .B1(_1613_),
    .B2(_1614_),
    .X(_1620_));
 sky130_fd_sc_hd__nand4_2 _5873_ (.A(_1613_),
    .B(_1614_),
    .C(net226),
    .D(net317),
    .Y(_1621_));
 sky130_fd_sc_hd__o22ai_4 _5874_ (.A1(_1498_),
    .A2(_1608_),
    .B1(_1609_),
    .B2(_1548_),
    .Y(_1622_));
 sky130_fd_sc_hd__nand3_4 _5875_ (.A(_1620_),
    .B(_1621_),
    .C(_1622_),
    .Y(_1623_));
 sky130_fd_sc_hd__a21bo_1 _5876_ (.A1(_1554_),
    .A2(_1557_),
    .B1_N(_1555_),
    .X(_1624_));
 sky130_fd_sc_hd__nand3_4 _5877_ (.A(_1619_),
    .B(_1623_),
    .C(_1624_),
    .Y(_1625_));
 sky130_fd_sc_hd__o32a_1 _5878_ (.A1(_0385_),
    .A2(_1415_),
    .A3(_1481_),
    .B1(_3441_),
    .B2(_1332_),
    .X(_1626_));
 sky130_fd_sc_hd__o22a_1 _5879_ (.A1(_1355_),
    .A2(_0385_),
    .B1(_1415_),
    .B2(_3134_),
    .X(_1627_));
 sky130_fd_sc_hd__o2bb2ai_4 _5880_ (.A1_N(_1619_),
    .A2_N(_1623_),
    .B1(_1626_),
    .B2(_1627_),
    .Y(_1628_));
 sky130_fd_sc_hd__nand2_4 _5881_ (.A(net392),
    .B(net190),
    .Y(_1630_));
 sky130_fd_sc_hd__nand2_2 _5882_ (.A(net366),
    .B(net201),
    .Y(_1631_));
 sky130_fd_sc_hd__nand2_2 _5883_ (.A(_1608_),
    .B(_1631_),
    .Y(_1632_));
 sky130_fd_sc_hd__nand4_4 _5884_ (.A(net378),
    .B(net370),
    .C(net202),
    .D(net195),
    .Y(_1633_));
 sky130_fd_sc_hd__o211ai_4 _5885_ (.A1(_3134_),
    .A2(_1393_),
    .B1(_1632_),
    .C1(_1633_),
    .Y(_1634_));
 sky130_fd_sc_hd__nand2_1 _5886_ (.A(net357),
    .B(net208),
    .Y(_1635_));
 sky130_fd_sc_hd__a21o_2 _5887_ (.A1(_1632_),
    .A2(_1633_),
    .B1(_1635_),
    .X(_1636_));
 sky130_fd_sc_hd__and3_1 _5888_ (.A(_1630_),
    .B(_1634_),
    .C(_1636_),
    .X(_1637_));
 sky130_fd_sc_hd__a21oi_4 _5889_ (.A1(_1634_),
    .A2(_1636_),
    .B1(_1630_),
    .Y(_1638_));
 sky130_fd_sc_hd__o2bb2ai_4 _5890_ (.A1_N(_1625_),
    .A2_N(_1628_),
    .B1(_1637_),
    .B2(_1638_),
    .Y(_1639_));
 sky130_fd_sc_hd__inv_4 _5891_ (.A(net192),
    .Y(_1641_));
 sky130_fd_sc_hd__buf_6 _5892_ (.A(_1641_),
    .X(_1642_));
 sky130_fd_sc_hd__buf_4 _5893_ (.A(_1642_),
    .X(_1643_));
 sky130_fd_sc_hd__o211ai_4 _5894_ (.A1(_1329_),
    .A2(_1643_),
    .B1(_1634_),
    .C1(_1636_),
    .Y(_1644_));
 sky130_fd_sc_hd__a22oi_1 _5895_ (.A1(net354),
    .A2(net208),
    .B1(_1632_),
    .B2(_1633_),
    .Y(_1645_));
 sky130_fd_sc_hd__nand4_1 _5896_ (.A(_1632_),
    .B(_1633_),
    .C(net354),
    .D(net208),
    .Y(_1646_));
 sky130_fd_sc_hd__nor2_1 _5897_ (.A(_3125_),
    .B(_1643_),
    .Y(_1647_));
 sky130_fd_sc_hd__nand3b_4 _5898_ (.A_N(_1645_),
    .B(_1646_),
    .C(_1647_),
    .Y(_1648_));
 sky130_fd_sc_hd__nand4_4 _5899_ (.A(_1625_),
    .B(_1628_),
    .C(_1644_),
    .D(_1648_),
    .Y(_1649_));
 sky130_fd_sc_hd__a21oi_4 _5900_ (.A1(_1571_),
    .A2(_1573_),
    .B1(_1574_),
    .Y(_1650_));
 sky130_fd_sc_hd__a21oi_4 _5901_ (.A1(_1639_),
    .A2(_1649_),
    .B1(_1650_),
    .Y(_1652_));
 sky130_fd_sc_hd__and3_2 _5902_ (.A(_1619_),
    .B(_1623_),
    .C(_1624_),
    .X(_1653_));
 sky130_fd_sc_hd__nand3_2 _5903_ (.A(_1628_),
    .B(_1644_),
    .C(_1648_),
    .Y(_1654_));
 sky130_fd_sc_hd__o211a_1 _5904_ (.A1(_1653_),
    .A2(_1654_),
    .B1(_1650_),
    .C1(_1639_),
    .X(_1655_));
 sky130_fd_sc_hd__a22oi_4 _5905_ (.A1(net235),
    .A2(net316),
    .B1(net306),
    .B2(net242),
    .Y(_1656_));
 sky130_fd_sc_hd__o21ai_1 _5906_ (.A1(_1530_),
    .A2(_1656_),
    .B1(_1526_),
    .Y(_1657_));
 sky130_fd_sc_hd__nand2_1 _5907_ (.A(net299),
    .B(net242),
    .Y(_1658_));
 sky130_fd_sc_hd__nand2_2 _5908_ (.A(_1533_),
    .B(_1658_),
    .Y(_1659_));
 sky130_fd_sc_hd__nand4_4 _5909_ (.A(net299),
    .B(net242),
    .C(net235),
    .D(net306),
    .Y(_1660_));
 sky130_fd_sc_hd__nand4_2 _5910_ (.A(_1659_),
    .B(net248),
    .C(net287),
    .D(_1660_),
    .Y(_1661_));
 sky130_fd_sc_hd__nand2_2 _5911_ (.A(_1657_),
    .B(_1661_),
    .Y(_1663_));
 sky130_fd_sc_hd__o2bb2a_2 _5912_ (.A1_N(_1660_),
    .A2_N(_1659_),
    .B1(_0509_),
    .B2(_1301_),
    .X(_1664_));
 sky130_fd_sc_hd__o22a_2 _5913_ (.A1(_3022_),
    .A2(_1129_),
    .B1(_1527_),
    .B2(_1528_),
    .X(_1665_));
 sky130_fd_sc_hd__nand2_4 _5914_ (.A(net300),
    .B(net234),
    .Y(_1666_));
 sky130_fd_sc_hd__o221ai_4 _5915_ (.A1(_3381_),
    .A2(_1129_),
    .B1(_1528_),
    .B2(_1666_),
    .C1(_1659_),
    .Y(_1667_));
 sky130_fd_sc_hd__nand2_1 _5916_ (.A(net287),
    .B(net248),
    .Y(_1668_));
 sky130_fd_sc_hd__a21o_1 _5917_ (.A1(_1660_),
    .A2(_1659_),
    .B1(_1668_),
    .X(_1669_));
 sky130_fd_sc_hd__o211ai_4 _5918_ (.A1(_1656_),
    .A2(_1665_),
    .B1(_1667_),
    .C1(_1669_),
    .Y(_1670_));
 sky130_fd_sc_hd__nand2_1 _5919_ (.A(_1563_),
    .B(_1572_),
    .Y(_1671_));
 sky130_fd_sc_hd__o2111ai_4 _5920_ (.A1(_1663_),
    .A2(_1664_),
    .B1(_1560_),
    .C1(_1670_),
    .D1(_1671_),
    .Y(_1672_));
 sky130_fd_sc_hd__o21ai_1 _5921_ (.A1(_1664_),
    .A2(_1663_),
    .B1(_1670_),
    .Y(_1674_));
 sky130_fd_sc_hd__a31o_1 _5922_ (.A1(_1551_),
    .A2(_1558_),
    .A3(_1559_),
    .B1(_1572_),
    .X(_1675_));
 sky130_fd_sc_hd__nand3_1 _5923_ (.A(_1563_),
    .B(_1674_),
    .C(_1675_),
    .Y(_1676_));
 sky130_fd_sc_hd__and4_1 _5924_ (.A(_1529_),
    .B(net247),
    .C(net299),
    .D(_1526_),
    .X(_1677_));
 sky130_fd_sc_hd__nand2_1 _5925_ (.A(_1536_),
    .B(_1525_),
    .Y(_1678_));
 sky130_fd_sc_hd__o2bb2ai_1 _5926_ (.A1_N(_1672_),
    .A2_N(_1676_),
    .B1(_1677_),
    .B2(_1678_),
    .Y(_1679_));
 sky130_fd_sc_hd__nand3b_1 _5927_ (.A_N(_1538_),
    .B(_1672_),
    .C(_1676_),
    .Y(_1680_));
 sky130_fd_sc_hd__nand2_2 _5928_ (.A(_1679_),
    .B(_1680_),
    .Y(_1681_));
 sky130_fd_sc_hd__o21bai_1 _5929_ (.A1(_1652_),
    .A2(_1655_),
    .B1_N(_1681_),
    .Y(_1682_));
 sky130_fd_sc_hd__a21o_1 _5930_ (.A1(_1591_),
    .A2(_1583_),
    .B1(_1578_),
    .X(_1683_));
 sky130_fd_sc_hd__a21o_1 _5931_ (.A1(_1639_),
    .A2(_1649_),
    .B1(_1650_),
    .X(_1685_));
 sky130_fd_sc_hd__o211ai_4 _5932_ (.A1(_1653_),
    .A2(_1654_),
    .B1(_1650_),
    .C1(_1639_),
    .Y(_1686_));
 sky130_fd_sc_hd__nand3_1 _5933_ (.A(_1685_),
    .B(_1686_),
    .C(_1681_),
    .Y(_1687_));
 sky130_fd_sc_hd__nand3_1 _5934_ (.A(_1682_),
    .B(_1683_),
    .C(_1687_),
    .Y(_1688_));
 sky130_fd_sc_hd__o21ai_1 _5935_ (.A1(_1652_),
    .A2(_1655_),
    .B1(_1681_),
    .Y(_1689_));
 sky130_fd_sc_hd__nand4_1 _5936_ (.A(_1685_),
    .B(_1686_),
    .C(_1679_),
    .D(_1680_),
    .Y(_1690_));
 sky130_fd_sc_hd__a21oi_1 _5937_ (.A1(_1591_),
    .A2(_1583_),
    .B1(_1578_),
    .Y(_1691_));
 sky130_fd_sc_hd__nand3_1 _5938_ (.A(_1689_),
    .B(_1690_),
    .C(_1691_),
    .Y(_1692_));
 sky130_fd_sc_hd__o21ai_1 _5939_ (.A1(_1490_),
    .A2(_1539_),
    .B1(_1541_),
    .Y(_1693_));
 sky130_fd_sc_hd__a21oi_2 _5940_ (.A1(_1688_),
    .A2(_1692_),
    .B1(_1693_),
    .Y(_1694_));
 sky130_fd_sc_hd__o211a_1 _5941_ (.A1(_1540_),
    .A2(_1543_),
    .B1(_1688_),
    .C1(_1692_),
    .X(_1696_));
 sky130_fd_sc_hd__nor2_1 _5942_ (.A(_1694_),
    .B(_1696_),
    .Y(_1697_));
 sky130_fd_sc_hd__xor2_1 _5943_ (.A(_1606_),
    .B(_1697_),
    .X(_1698_));
 sky130_fd_sc_hd__xnor2_1 _5944_ (.A(_1605_),
    .B(_1698_),
    .Y(_0104_));
 sky130_fd_sc_hd__nand2_1 _5945_ (.A(net287),
    .B(net242),
    .Y(_1699_));
 sky130_fd_sc_hd__nand2_1 _5946_ (.A(_1666_),
    .B(_1699_),
    .Y(_1700_));
 sky130_fd_sc_hd__nand4_2 _5947_ (.A(net299),
    .B(net287),
    .C(net242),
    .D(net235),
    .Y(_1701_));
 sky130_fd_sc_hd__a22oi_1 _5948_ (.A1(net274),
    .A2(net248),
    .B1(_1700_),
    .B2(_1701_),
    .Y(_1702_));
 sky130_fd_sc_hd__and4_1 _5949_ (.A(_1700_),
    .B(_1701_),
    .C(net274),
    .D(net248),
    .X(_1703_));
 sky130_fd_sc_hd__a22oi_2 _5950_ (.A1(_1533_),
    .A2(_1658_),
    .B1(_1660_),
    .B2(_1668_),
    .Y(_1704_));
 sky130_fd_sc_hd__o21bai_1 _5951_ (.A1(_1702_),
    .A2(_1703_),
    .B1_N(_1704_),
    .Y(_1706_));
 sky130_fd_sc_hd__a22o_1 _5952_ (.A1(net274),
    .A2(net248),
    .B1(_1700_),
    .B2(_1701_),
    .X(_1707_));
 sky130_fd_sc_hd__nand2_1 _5953_ (.A(net287),
    .B(net235),
    .Y(_1708_));
 sky130_fd_sc_hd__o2111ai_1 _5954_ (.A1(_1658_),
    .A2(_1708_),
    .B1(net274),
    .C1(net248),
    .D1(_1700_),
    .Y(_1709_));
 sky130_fd_sc_hd__nand3_1 _5955_ (.A(_1707_),
    .B(_1709_),
    .C(_1704_),
    .Y(_1710_));
 sky130_fd_sc_hd__nand2_2 _5956_ (.A(_1706_),
    .B(_1710_),
    .Y(_1711_));
 sky130_fd_sc_hd__a21oi_2 _5957_ (.A1(_1623_),
    .A2(_1625_),
    .B1(_1711_),
    .Y(_1712_));
 sky130_fd_sc_hd__o2bb2a_1 _5958_ (.A1_N(_1613_),
    .A2_N(_1614_),
    .B1(_1332_),
    .B2(net96),
    .X(_1713_));
 sky130_fd_sc_hd__nand2_1 _5959_ (.A(_1622_),
    .B(_1621_),
    .Y(_1714_));
 sky130_fd_sc_hd__o211a_2 _5960_ (.A1(_1713_),
    .A2(_1714_),
    .B1(_1625_),
    .C1(_1711_),
    .X(_1715_));
 sky130_fd_sc_hd__o22ai_2 _5961_ (.A1(_1664_),
    .A2(_1663_),
    .B1(_1712_),
    .B2(_1715_),
    .Y(_1717_));
 sky130_fd_sc_hd__a211o_1 _5962_ (.A1(_1667_),
    .A2(_1669_),
    .B1(_1656_),
    .C1(_1665_),
    .X(_1718_));
 sky130_fd_sc_hd__a21o_1 _5963_ (.A1(_1623_),
    .A2(_1625_),
    .B1(_1711_),
    .X(_1719_));
 sky130_fd_sc_hd__o211ai_4 _5964_ (.A1(_1713_),
    .A2(_1714_),
    .B1(_1625_),
    .C1(_1711_),
    .Y(_1720_));
 sky130_fd_sc_hd__nand3b_1 _5965_ (.A_N(_1718_),
    .B(_1719_),
    .C(_1720_),
    .Y(_1721_));
 sky130_fd_sc_hd__nand2_2 _5966_ (.A(_1717_),
    .B(_1721_),
    .Y(_1722_));
 sky130_fd_sc_hd__nand4_4 _5967_ (.A(net366),
    .B(net353),
    .C(net201),
    .D(net195),
    .Y(_1723_));
 sky130_fd_sc_hd__nand2_2 _5968_ (.A(net377),
    .B(net195),
    .Y(_1724_));
 sky130_fd_sc_hd__nand2_1 _5969_ (.A(net353),
    .B(net201),
    .Y(_1725_));
 sky130_fd_sc_hd__nand2_2 _5970_ (.A(_1724_),
    .B(_1725_),
    .Y(_1726_));
 sky130_fd_sc_hd__nand2_2 _5971_ (.A(net342),
    .B(net208),
    .Y(_1728_));
 sky130_fd_sc_hd__a21oi_2 _5972_ (.A1(_1723_),
    .A2(_1726_),
    .B1(_1728_),
    .Y(_1729_));
 sky130_fd_sc_hd__a22oi_4 _5973_ (.A1(net354),
    .A2(net201),
    .B1(net195),
    .B2(net366),
    .Y(_1730_));
 sky130_fd_sc_hd__nand2_2 _5974_ (.A(_1728_),
    .B(_1723_),
    .Y(_1731_));
 sky130_fd_sc_hd__nand2_2 _5975_ (.A(net378),
    .B(net182),
    .Y(_1732_));
 sky130_fd_sc_hd__nand2_1 _5976_ (.A(net392),
    .B(net182),
    .Y(_1733_));
 sky130_fd_sc_hd__nand2_1 _5977_ (.A(net378),
    .B(net190),
    .Y(_1734_));
 sky130_fd_sc_hd__nand2_1 _5978_ (.A(_1733_),
    .B(_1734_),
    .Y(_1735_));
 sky130_fd_sc_hd__o21ai_4 _5979_ (.A1(_1630_),
    .A2(_1732_),
    .B1(_1735_),
    .Y(_1736_));
 sky130_fd_sc_hd__o21ai_2 _5980_ (.A1(_1730_),
    .A2(_1731_),
    .B1(_1736_),
    .Y(_1737_));
 sky130_fd_sc_hd__o2bb2ai_1 _5981_ (.A1_N(_1723_),
    .A2_N(_1726_),
    .B1(_0385_),
    .B2(_1393_),
    .Y(_1739_));
 sky130_fd_sc_hd__o21a_1 _5982_ (.A1(_1630_),
    .A2(_1732_),
    .B1(_1735_),
    .X(_1740_));
 sky130_fd_sc_hd__nand4_1 _5983_ (.A(_1726_),
    .B(net208),
    .C(net340),
    .D(_1723_),
    .Y(_1741_));
 sky130_fd_sc_hd__nand3_2 _5984_ (.A(_1739_),
    .B(_1740_),
    .C(_1741_),
    .Y(_1742_));
 sky130_fd_sc_hd__o21ai_2 _5985_ (.A1(_1729_),
    .A2(_1737_),
    .B1(_1742_),
    .Y(_1743_));
 sky130_fd_sc_hd__nand2_2 _5986_ (.A(_1648_),
    .B(_1743_),
    .Y(_1744_));
 sky130_fd_sc_hd__o211ai_4 _5987_ (.A1(_1729_),
    .A2(_1737_),
    .B1(_1742_),
    .C1(_1638_),
    .Y(_1745_));
 sky130_fd_sc_hd__nand4_4 _5988_ (.A(net220),
    .B(net215),
    .C(net330),
    .D(net318),
    .Y(_1746_));
 sky130_fd_sc_hd__nand2_1 _5989_ (.A(net214),
    .B(net339),
    .Y(_1747_));
 sky130_fd_sc_hd__nand2_1 _5990_ (.A(net220),
    .B(net318),
    .Y(_1748_));
 sky130_fd_sc_hd__nand2_4 _5991_ (.A(_1747_),
    .B(_1748_),
    .Y(_1750_));
 sky130_fd_sc_hd__nand2_2 _5992_ (.A(net226),
    .B(net308),
    .Y(_1751_));
 sky130_fd_sc_hd__a21oi_4 _5993_ (.A1(_1746_),
    .A2(_1750_),
    .B1(_1751_),
    .Y(_1752_));
 sky130_fd_sc_hd__a22o_1 _5994_ (.A1(_1608_),
    .A2(_1631_),
    .B1(_1633_),
    .B2(_1635_),
    .X(_1753_));
 sky130_fd_sc_hd__o211ai_1 _5995_ (.A1(_1366_),
    .A2(_2848_),
    .B1(_1746_),
    .C1(_1750_),
    .Y(_1754_));
 sky130_fd_sc_hd__nand2_2 _5996_ (.A(_1753_),
    .B(_1754_),
    .Y(_1755_));
 sky130_fd_sc_hd__o2bb2ai_1 _5997_ (.A1_N(_1746_),
    .A2_N(_1750_),
    .B1(_1366_),
    .B2(_2848_),
    .Y(_1756_));
 sky130_fd_sc_hd__nand4_1 _5998_ (.A(_1750_),
    .B(net307),
    .C(net226),
    .D(_1746_),
    .Y(_1757_));
 sky130_fd_sc_hd__a22oi_1 _5999_ (.A1(_1608_),
    .A2(_1631_),
    .B1(_1633_),
    .B2(_1635_),
    .Y(_1758_));
 sky130_fd_sc_hd__nand3_1 _6000_ (.A(_1756_),
    .B(_1757_),
    .C(_1758_),
    .Y(_1759_));
 sky130_fd_sc_hd__buf_2 _6001_ (.A(_1759_),
    .X(_1761_));
 sky130_fd_sc_hd__o21a_1 _6002_ (.A1(_2965_),
    .A2(_1367_),
    .B1(_1612_),
    .X(_1762_));
 sky130_fd_sc_hd__o32a_2 _6003_ (.A1(_1415_),
    .A2(_3441_),
    .A3(_1552_),
    .B1(_1616_),
    .B2(_1762_),
    .X(_1763_));
 sky130_fd_sc_hd__o211a_1 _6004_ (.A1(_1752_),
    .A2(_1755_),
    .B1(_1761_),
    .C1(_1763_),
    .X(_1764_));
 sky130_fd_sc_hd__nand2_2 _6005_ (.A(net219),
    .B(net318),
    .Y(_1765_));
 sky130_fd_sc_hd__o21ai_4 _6006_ (.A1(_1612_),
    .A2(_1765_),
    .B1(_1751_),
    .Y(_1766_));
 sky130_fd_sc_hd__a22oi_4 _6007_ (.A1(net215),
    .A2(net329),
    .B1(net317),
    .B2(net221),
    .Y(_1767_));
 sky130_fd_sc_hd__a21o_1 _6008_ (.A1(_1746_),
    .A2(_1750_),
    .B1(_1751_),
    .X(_1768_));
 sky130_fd_sc_hd__o211ai_4 _6009_ (.A1(_1766_),
    .A2(_1767_),
    .B1(_1753_),
    .C1(_1768_),
    .Y(_1769_));
 sky130_fd_sc_hd__a21oi_1 _6010_ (.A1(_1761_),
    .A2(_1769_),
    .B1(_1763_),
    .Y(_1770_));
 sky130_fd_sc_hd__o2bb2ai_1 _6011_ (.A1_N(_1744_),
    .A2_N(_1745_),
    .B1(_1764_),
    .B2(_1770_),
    .Y(_1772_));
 sky130_fd_sc_hd__o2111ai_1 _6012_ (.A1(_1616_),
    .A2(_1762_),
    .B1(_1614_),
    .C1(_1761_),
    .D1(_1769_),
    .Y(_1773_));
 sky130_fd_sc_hd__o21ai_2 _6013_ (.A1(_1752_),
    .A2(_1755_),
    .B1(_1759_),
    .Y(_1774_));
 sky130_fd_sc_hd__o21ai_2 _6014_ (.A1(_1616_),
    .A2(_1762_),
    .B1(_1614_),
    .Y(_1775_));
 sky130_fd_sc_hd__nand2_1 _6015_ (.A(_1774_),
    .B(_1775_),
    .Y(_1776_));
 sky130_fd_sc_hd__nand4_1 _6016_ (.A(_1744_),
    .B(_1745_),
    .C(_1773_),
    .D(_1776_),
    .Y(_1777_));
 sky130_fd_sc_hd__o211ai_2 _6017_ (.A1(_1653_),
    .A2(_1654_),
    .B1(_1772_),
    .C1(_1777_),
    .Y(_1778_));
 sky130_fd_sc_hd__nand2_1 _6018_ (.A(_1644_),
    .B(_1648_),
    .Y(_1779_));
 sky130_fd_sc_hd__a21oi_1 _6019_ (.A1(_1619_),
    .A2(_1623_),
    .B1(_1624_),
    .Y(_1780_));
 sky130_fd_sc_hd__nor3_1 _6020_ (.A(_1779_),
    .B(_1780_),
    .C(_1653_),
    .Y(_1781_));
 sky130_fd_sc_hd__o211a_1 _6021_ (.A1(_1752_),
    .A2(_1755_),
    .B1(_1761_),
    .C1(_1775_),
    .X(_1783_));
 sky130_fd_sc_hd__a21oi_2 _6022_ (.A1(_1761_),
    .A2(_1769_),
    .B1(_1775_),
    .Y(_1784_));
 sky130_fd_sc_hd__o2bb2ai_1 _6023_ (.A1_N(_1744_),
    .A2_N(_1745_),
    .B1(_1783_),
    .B2(_1784_),
    .Y(_1785_));
 sky130_fd_sc_hd__o211ai_2 _6024_ (.A1(_1752_),
    .A2(_1755_),
    .B1(_1761_),
    .C1(_1775_),
    .Y(_1786_));
 sky130_fd_sc_hd__nand2_1 _6025_ (.A(_1763_),
    .B(_1774_),
    .Y(_1787_));
 sky130_fd_sc_hd__nand4_1 _6026_ (.A(_1744_),
    .B(_1745_),
    .C(_1786_),
    .D(_1787_),
    .Y(_1788_));
 sky130_fd_sc_hd__nand3_1 _6027_ (.A(_1781_),
    .B(_1785_),
    .C(_1788_),
    .Y(_1789_));
 sky130_fd_sc_hd__nand3_1 _6028_ (.A(_1722_),
    .B(_1778_),
    .C(_1789_),
    .Y(_1790_));
 sky130_fd_sc_hd__a21oi_1 _6029_ (.A1(_1719_),
    .A2(_1720_),
    .B1(_1718_),
    .Y(_1791_));
 sky130_fd_sc_hd__a22o_1 _6030_ (.A1(net287),
    .A2(net248),
    .B1(_1660_),
    .B2(_1659_),
    .X(_1792_));
 sky130_fd_sc_hd__nand2_1 _6031_ (.A(_1792_),
    .B(_1661_),
    .Y(_1794_));
 sky130_fd_sc_hd__o311a_1 _6032_ (.A1(_1656_),
    .A2(_1665_),
    .A3(_1794_),
    .B1(_1719_),
    .C1(_1720_),
    .X(_1795_));
 sky130_fd_sc_hd__nand2_1 _6033_ (.A(_1778_),
    .B(_1789_),
    .Y(_1796_));
 sky130_fd_sc_hd__o21ai_1 _6034_ (.A1(_1791_),
    .A2(_1795_),
    .B1(_1796_),
    .Y(_1797_));
 sky130_fd_sc_hd__o2111ai_4 _6035_ (.A1(_1681_),
    .A2(_1652_),
    .B1(_1686_),
    .C1(_1790_),
    .D1(_1797_),
    .Y(_1798_));
 sky130_fd_sc_hd__o21ai_1 _6036_ (.A1(_1652_),
    .A2(_1681_),
    .B1(_1686_),
    .Y(_1799_));
 sky130_fd_sc_hd__nand4_1 _6037_ (.A(_1717_),
    .B(_1721_),
    .C(_1778_),
    .D(_1789_),
    .Y(_1800_));
 sky130_fd_sc_hd__nand2_1 _6038_ (.A(_1722_),
    .B(_1796_),
    .Y(_1801_));
 sky130_fd_sc_hd__nand3_2 _6039_ (.A(_1799_),
    .B(_1800_),
    .C(_1801_),
    .Y(_1802_));
 sky130_fd_sc_hd__nand2_1 _6040_ (.A(_1798_),
    .B(_1802_),
    .Y(_1803_));
 sky130_fd_sc_hd__a31o_1 _6041_ (.A1(_1563_),
    .A2(_1674_),
    .A3(_1675_),
    .B1(_1538_),
    .X(_1805_));
 sky130_fd_sc_hd__nand2_1 _6042_ (.A(_1672_),
    .B(_1805_),
    .Y(_1806_));
 sky130_fd_sc_hd__nand2_1 _6043_ (.A(_1803_),
    .B(_1806_),
    .Y(_1807_));
 sky130_fd_sc_hd__nand4_1 _6044_ (.A(_1672_),
    .B(_1798_),
    .C(_1802_),
    .D(_1805_),
    .Y(_1808_));
 sky130_fd_sc_hd__nand2_2 _6045_ (.A(_1807_),
    .B(_1808_),
    .Y(_1809_));
 sky130_fd_sc_hd__a32o_2 _6046_ (.A1(_1689_),
    .A2(_1690_),
    .A3(_1691_),
    .B1(_1688_),
    .B2(_1693_),
    .X(_1810_));
 sky130_fd_sc_hd__and2_1 _6047_ (.A(_1809_),
    .B(_1810_),
    .X(_1811_));
 sky130_fd_sc_hd__nor2_1 _6048_ (.A(_1810_),
    .B(_1809_),
    .Y(_1812_));
 sky130_fd_sc_hd__or2_1 _6049_ (.A(_1811_),
    .B(_1812_),
    .X(_1813_));
 sky130_fd_sc_hd__or2_1 _6050_ (.A(_1694_),
    .B(_1696_),
    .X(_1814_));
 sky130_fd_sc_hd__a21bo_1 _6051_ (.A1(_1594_),
    .A2(_1599_),
    .B1_N(_1589_),
    .X(_1816_));
 sky130_fd_sc_hd__a21o_1 _6052_ (.A1(_1598_),
    .A2(_1600_),
    .B1(_1602_),
    .X(_1817_));
 sky130_fd_sc_hd__nand2_1 _6053_ (.A(_1522_),
    .B(_1604_),
    .Y(_1818_));
 sky130_fd_sc_hd__o211ai_2 _6054_ (.A1(_1816_),
    .A2(_1697_),
    .B1(_1817_),
    .C1(_1818_),
    .Y(_1819_));
 sky130_fd_sc_hd__o21ai_1 _6055_ (.A1(_1606_),
    .A2(_1814_),
    .B1(_1819_),
    .Y(_1820_));
 sky130_fd_sc_hd__xnor2_1 _6056_ (.A(_1813_),
    .B(_1820_),
    .Y(_0087_));
 sky130_fd_sc_hd__nand2_1 _6057_ (.A(net209),
    .B(net330),
    .Y(_1821_));
 sky130_fd_sc_hd__nand2_2 _6058_ (.A(_1765_),
    .B(_1821_),
    .Y(_1822_));
 sky130_fd_sc_hd__nand4_4 _6059_ (.A(net209),
    .B(net218),
    .C(net330),
    .D(net318),
    .Y(_1823_));
 sky130_fd_sc_hd__o2bb2ai_4 _6060_ (.A1_N(_1822_),
    .A2_N(_1823_),
    .B1(_1355_),
    .B2(_2783_),
    .Y(_1824_));
 sky130_fd_sc_hd__nand4_4 _6061_ (.A(_1822_),
    .B(_1823_),
    .C(net225),
    .D(net308),
    .Y(_1826_));
 sky130_fd_sc_hd__nand2_2 _6062_ (.A(net353),
    .B(net195),
    .Y(_1827_));
 sky130_fd_sc_hd__o22ai_4 _6063_ (.A1(_1631_),
    .A2(_1827_),
    .B1(_1728_),
    .B2(_1730_),
    .Y(_1828_));
 sky130_fd_sc_hd__and3_1 _6064_ (.A(_1824_),
    .B(_1826_),
    .C(_1828_),
    .X(_1829_));
 sky130_fd_sc_hd__clkbuf_4 _6065_ (.A(_1829_),
    .X(_1830_));
 sky130_fd_sc_hd__a21o_1 _6066_ (.A1(_1824_),
    .A2(_1826_),
    .B1(_1828_),
    .X(_1831_));
 sky130_fd_sc_hd__o32a_1 _6067_ (.A1(_1367_),
    .A2(_1782_),
    .A3(_1612_),
    .B1(_1751_),
    .B2(_1767_),
    .X(_1832_));
 sky130_fd_sc_hd__inv_2 _6068_ (.A(_1832_),
    .Y(_1833_));
 sky130_fd_sc_hd__nand2_2 _6069_ (.A(_1831_),
    .B(_1833_),
    .Y(_1834_));
 sky130_fd_sc_hd__a21oi_2 _6070_ (.A1(_1824_),
    .A2(_1826_),
    .B1(_1828_),
    .Y(_1835_));
 sky130_fd_sc_hd__o21bai_4 _6071_ (.A1(_1835_),
    .A2(_1830_),
    .B1_N(_1833_),
    .Y(_1837_));
 sky130_fd_sc_hd__o21ai_2 _6072_ (.A1(_1830_),
    .A2(_1834_),
    .B1(_1837_),
    .Y(_1838_));
 sky130_fd_sc_hd__nand2_1 _6073_ (.A(net366),
    .B(net190),
    .Y(_1839_));
 sky130_fd_sc_hd__nand2_4 _6074_ (.A(_1827_),
    .B(_1839_),
    .Y(_1840_));
 sky130_fd_sc_hd__nand4_1 _6075_ (.A(net366),
    .B(net353),
    .C(net195),
    .D(net190),
    .Y(_1841_));
 sky130_fd_sc_hd__a22o_1 _6076_ (.A1(net340),
    .A2(net201),
    .B1(_1840_),
    .B2(_1841_),
    .X(_1842_));
 sky130_fd_sc_hd__o211ai_1 _6077_ (.A1(net190),
    .A2(_1732_),
    .B1(net178),
    .C1(net392),
    .Y(_1843_));
 sky130_fd_sc_hd__nand2_1 _6078_ (.A(net392),
    .B(net178),
    .Y(_1844_));
 sky130_fd_sc_hd__nand4_2 _6079_ (.A(_1630_),
    .B(_1844_),
    .C(net378),
    .D(net182),
    .Y(_1845_));
 sky130_fd_sc_hd__nand2_1 _6080_ (.A(_1843_),
    .B(_1845_),
    .Y(_1846_));
 sky130_fd_sc_hd__nand2_4 _6081_ (.A(net353),
    .B(net190),
    .Y(_1848_));
 sky130_fd_sc_hd__o2111ai_4 _6082_ (.A1(_1724_),
    .A2(_1848_),
    .B1(net340),
    .C1(net207),
    .D1(_1840_),
    .Y(_1849_));
 sky130_fd_sc_hd__nand3_4 _6083_ (.A(_1842_),
    .B(_1846_),
    .C(_1849_),
    .Y(_1850_));
 sky130_fd_sc_hd__o21ai_1 _6084_ (.A1(net190),
    .A2(_1732_),
    .B1(net178),
    .Y(_1851_));
 sky130_fd_sc_hd__nand2_1 _6085_ (.A(net340),
    .B(net207),
    .Y(_1852_));
 sky130_fd_sc_hd__o211ai_2 _6086_ (.A1(_1724_),
    .A2(_1848_),
    .B1(_1840_),
    .C1(_1852_),
    .Y(_1853_));
 sky130_fd_sc_hd__a21o_1 _6087_ (.A1(_1840_),
    .A2(_1841_),
    .B1(_1852_),
    .X(_1854_));
 sky130_fd_sc_hd__o2111ai_4 _6088_ (.A1(_3125_),
    .A2(_1851_),
    .B1(_1845_),
    .C1(_1853_),
    .D1(_1854_),
    .Y(_1855_));
 sky130_fd_sc_hd__nand3b_4 _6089_ (.A_N(_1742_),
    .B(_1850_),
    .C(_1855_),
    .Y(_1856_));
 sky130_fd_sc_hd__nand2_1 _6090_ (.A(_1739_),
    .B(_1741_),
    .Y(_1857_));
 sky130_fd_sc_hd__o2bb2ai_4 _6091_ (.A1_N(_1850_),
    .A2_N(_1855_),
    .B1(_1857_),
    .B2(_1736_),
    .Y(_1859_));
 sky130_fd_sc_hd__nand2_1 _6092_ (.A(_1856_),
    .B(_1859_),
    .Y(_1860_));
 sky130_fd_sc_hd__nand2_1 _6093_ (.A(_1838_),
    .B(_1860_),
    .Y(_1861_));
 sky130_fd_sc_hd__o2bb2ai_1 _6094_ (.A1_N(_1648_),
    .A2_N(_1743_),
    .B1(_1763_),
    .B2(_1774_),
    .Y(_1862_));
 sky130_fd_sc_hd__o21ai_2 _6095_ (.A1(_1784_),
    .A2(_1862_),
    .B1(_1745_),
    .Y(_1863_));
 sky130_fd_sc_hd__o2111ai_4 _6096_ (.A1(_1830_),
    .A2(_1834_),
    .B1(_1856_),
    .C1(_1859_),
    .D1(_1837_),
    .Y(_1864_));
 sky130_fd_sc_hd__nand3_4 _6097_ (.A(_1861_),
    .B(_1863_),
    .C(_1864_),
    .Y(_1865_));
 sky130_fd_sc_hd__o22a_1 _6098_ (.A1(_1648_),
    .A2(_1743_),
    .B1(_1784_),
    .B2(_1862_),
    .X(_1866_));
 sky130_fd_sc_hd__nand3_1 _6099_ (.A(_1838_),
    .B(_1856_),
    .C(_1859_),
    .Y(_1867_));
 sky130_fd_sc_hd__o211ai_2 _6100_ (.A1(_1834_),
    .A2(_1830_),
    .B1(_1837_),
    .C1(_1860_),
    .Y(_1868_));
 sky130_fd_sc_hd__nand3_4 _6101_ (.A(_1866_),
    .B(_1867_),
    .C(_1868_),
    .Y(_1870_));
 sky130_fd_sc_hd__a2bb2o_2 _6102_ (.A1_N(_1752_),
    .A2_N(_1755_),
    .B1(_1759_),
    .B2(_1763_),
    .X(_1871_));
 sky130_fd_sc_hd__a22oi_4 _6103_ (.A1(net287),
    .A2(net242),
    .B1(net234),
    .B2(net300),
    .Y(_1872_));
 sky130_fd_sc_hd__nand2_1 _6104_ (.A(net274),
    .B(net249),
    .Y(_1873_));
 sky130_fd_sc_hd__o21a_1 _6105_ (.A1(_1666_),
    .A2(_1699_),
    .B1(_1873_),
    .X(_1874_));
 sky130_fd_sc_hd__nand2_2 _6106_ (.A(net288),
    .B(net229),
    .Y(_1875_));
 sky130_fd_sc_hd__a22o_1 _6107_ (.A1(net288),
    .A2(net234),
    .B1(net227),
    .B2(net300),
    .X(_1876_));
 sky130_fd_sc_hd__nand2_1 _6108_ (.A(net274),
    .B(net241),
    .Y(_1877_));
 sky130_fd_sc_hd__o211ai_2 _6109_ (.A1(_1666_),
    .A2(_1875_),
    .B1(_1876_),
    .C1(_1877_),
    .Y(_1878_));
 sky130_fd_sc_hd__nand2_1 _6110_ (.A(net300),
    .B(net228),
    .Y(_1879_));
 sky130_fd_sc_hd__o2bb2ai_1 _6111_ (.A1_N(_1708_),
    .A2_N(_1879_),
    .B1(_1875_),
    .B2(_1666_),
    .Y(_1881_));
 sky130_fd_sc_hd__nand3_1 _6112_ (.A(_1881_),
    .B(net241),
    .C(net274),
    .Y(_1882_));
 sky130_fd_sc_hd__o211ai_4 _6113_ (.A1(_1872_),
    .A2(_1874_),
    .B1(_1878_),
    .C1(_1882_),
    .Y(_1883_));
 sky130_fd_sc_hd__nand2_1 _6114_ (.A(_1877_),
    .B(_1881_),
    .Y(_1884_));
 sky130_fd_sc_hd__o2111ai_1 _6115_ (.A1(_1666_),
    .A2(_1875_),
    .B1(net274),
    .C1(net241),
    .D1(_1876_),
    .Y(_1885_));
 sky130_fd_sc_hd__o21ai_1 _6116_ (.A1(_1873_),
    .A2(_1872_),
    .B1(_1701_),
    .Y(_1886_));
 sky130_fd_sc_hd__nand3_2 _6117_ (.A(_1884_),
    .B(_1885_),
    .C(_1886_),
    .Y(_1887_));
 sky130_fd_sc_hd__o211ai_2 _6118_ (.A1(_3176_),
    .A2(_1301_),
    .B1(_1883_),
    .C1(_1887_),
    .Y(_1888_));
 sky130_fd_sc_hd__nand2_1 _6119_ (.A(net261),
    .B(net248),
    .Y(_1889_));
 sky130_fd_sc_hd__a21o_1 _6120_ (.A1(_1883_),
    .A2(_1887_),
    .B1(_1889_),
    .X(_1890_));
 sky130_fd_sc_hd__nand3_2 _6121_ (.A(_1871_),
    .B(_1888_),
    .C(_1890_),
    .Y(_1892_));
 sky130_fd_sc_hd__a22o_1 _6122_ (.A1(net261),
    .A2(net249),
    .B1(_1883_),
    .B2(_1887_),
    .X(_1893_));
 sky130_fd_sc_hd__nand4_1 _6123_ (.A(_1883_),
    .B(_1887_),
    .C(net261),
    .D(net249),
    .Y(_1894_));
 sky130_fd_sc_hd__a2bb2oi_2 _6124_ (.A1_N(_1752_),
    .A2_N(_1755_),
    .B1(_1761_),
    .B2(_1763_),
    .Y(_1895_));
 sky130_fd_sc_hd__nand3_1 _6125_ (.A(_1893_),
    .B(_1894_),
    .C(_1895_),
    .Y(_1896_));
 sky130_fd_sc_hd__and3_1 _6126_ (.A(_1707_),
    .B(_1709_),
    .C(_1704_),
    .X(_1897_));
 sky130_fd_sc_hd__a21oi_1 _6127_ (.A1(_1892_),
    .A2(_1896_),
    .B1(_1897_),
    .Y(_1898_));
 sky130_fd_sc_hd__nand3_1 _6128_ (.A(_1892_),
    .B(_1896_),
    .C(_1897_),
    .Y(_1899_));
 sky130_fd_sc_hd__inv_2 _6129_ (.A(_1899_),
    .Y(_1900_));
 sky130_fd_sc_hd__o2bb2ai_2 _6130_ (.A1_N(_1865_),
    .A2_N(_1870_),
    .B1(_1898_),
    .B2(_1900_),
    .Y(_1901_));
 sky130_fd_sc_hd__and3_1 _6131_ (.A(_1893_),
    .B(_1894_),
    .C(_1895_),
    .X(_1903_));
 sky130_fd_sc_hd__a31o_1 _6132_ (.A1(_1871_),
    .A2(_1888_),
    .A3(_1890_),
    .B1(_1710_),
    .X(_1904_));
 sky130_fd_sc_hd__a21o_1 _6133_ (.A1(_1892_),
    .A2(_1896_),
    .B1(_1897_),
    .X(_1905_));
 sky130_fd_sc_hd__o2111ai_4 _6134_ (.A1(_1903_),
    .A2(_1904_),
    .B1(_1905_),
    .C1(_1865_),
    .D1(_1870_),
    .Y(_1906_));
 sky130_fd_sc_hd__inv_2 _6135_ (.A(_1785_),
    .Y(_1907_));
 sky130_fd_sc_hd__a41o_1 _6136_ (.A1(_1744_),
    .A2(_1745_),
    .A3(_1786_),
    .A4(_1787_),
    .B1(_1649_),
    .X(_1908_));
 sky130_fd_sc_hd__o211a_1 _6137_ (.A1(_1653_),
    .A2(_1654_),
    .B1(_1772_),
    .C1(_1777_),
    .X(_1909_));
 sky130_fd_sc_hd__o22ai_4 _6138_ (.A1(_1907_),
    .A2(_1908_),
    .B1(_1909_),
    .B2(_1722_),
    .Y(_1910_));
 sky130_fd_sc_hd__a21o_1 _6139_ (.A1(_1901_),
    .A2(_1906_),
    .B1(_1910_),
    .X(_1911_));
 sky130_fd_sc_hd__nand3_1 _6140_ (.A(_1901_),
    .B(_1910_),
    .C(_1906_),
    .Y(_1912_));
 sky130_fd_sc_hd__a41o_1 _6141_ (.A1(_1792_),
    .A2(_1661_),
    .A3(_1720_),
    .A4(_1657_),
    .B1(_1712_),
    .X(_1914_));
 sky130_fd_sc_hd__nand3_2 _6142_ (.A(_1911_),
    .B(_1912_),
    .C(_1914_),
    .Y(_1915_));
 sky130_fd_sc_hd__o31a_1 _6143_ (.A1(_1656_),
    .A2(_1665_),
    .A3(_1794_),
    .B1(_1719_),
    .X(_1916_));
 sky130_fd_sc_hd__a21oi_2 _6144_ (.A1(_1901_),
    .A2(_1906_),
    .B1(_1910_),
    .Y(_1917_));
 sky130_fd_sc_hd__and3_1 _6145_ (.A(_1901_),
    .B(_1910_),
    .C(_1906_),
    .X(_1918_));
 sky130_fd_sc_hd__o22ai_4 _6146_ (.A1(_1715_),
    .A2(_1916_),
    .B1(_1917_),
    .B2(_1918_),
    .Y(_1919_));
 sky130_fd_sc_hd__nand2_1 _6147_ (.A(_1798_),
    .B(_1806_),
    .Y(_1920_));
 sky130_fd_sc_hd__nand2_2 _6148_ (.A(_1802_),
    .B(_1920_),
    .Y(_1921_));
 sky130_fd_sc_hd__a21oi_1 _6149_ (.A1(_1915_),
    .A2(_1919_),
    .B1(_1921_),
    .Y(_1922_));
 sky130_fd_sc_hd__and3_1 _6150_ (.A(_1919_),
    .B(_1921_),
    .C(_1915_),
    .X(_1923_));
 sky130_fd_sc_hd__nor2_1 _6151_ (.A(_1922_),
    .B(_1923_),
    .Y(_1925_));
 sky130_fd_sc_hd__or2_1 _6152_ (.A(_1810_),
    .B(_1809_),
    .X(_1926_));
 sky130_fd_sc_hd__a21oi_1 _6153_ (.A1(_1820_),
    .A2(_1926_),
    .B1(_1811_),
    .Y(_1927_));
 sky130_fd_sc_hd__xnor2_1 _6154_ (.A(_1925_),
    .B(_1927_),
    .Y(_0088_));
 sky130_fd_sc_hd__o2bb2a_2 _6155_ (.A1_N(_1850_),
    .A2_N(_1855_),
    .B1(_1857_),
    .B2(_1736_),
    .X(_1928_));
 sky130_fd_sc_hd__nand4_4 _6156_ (.A(_1726_),
    .B(_1731_),
    .C(_1824_),
    .D(_1826_),
    .Y(_1929_));
 sky130_fd_sc_hd__nand4_4 _6157_ (.A(_1750_),
    .B(_1766_),
    .C(_1831_),
    .D(_1929_),
    .Y(_1930_));
 sky130_fd_sc_hd__a21boi_1 _6158_ (.A1(_1837_),
    .A2(_1930_),
    .B1_N(_1856_),
    .Y(_1931_));
 sky130_fd_sc_hd__and2_1 _6159_ (.A(net340),
    .B(net201),
    .X(_1932_));
 sky130_fd_sc_hd__a21boi_4 _6160_ (.A1(_1840_),
    .A2(_1932_),
    .B1_N(_1841_),
    .Y(_1933_));
 sky130_fd_sc_hd__nand2_2 _6161_ (.A(net224),
    .B(net308),
    .Y(_1935_));
 sky130_fd_sc_hd__nand2_4 _6162_ (.A(net301),
    .B(net218),
    .Y(_1936_));
 sky130_fd_sc_hd__nand2_1 _6163_ (.A(net218),
    .B(net308),
    .Y(_1937_));
 sky130_fd_sc_hd__nand2_1 _6164_ (.A(net301),
    .B(net224),
    .Y(_1938_));
 sky130_fd_sc_hd__nand2_2 _6165_ (.A(_1937_),
    .B(_1938_),
    .Y(_1939_));
 sky130_fd_sc_hd__o2111ai_4 _6166_ (.A1(_1935_),
    .A2(_1936_),
    .B1(net287),
    .C1(net229),
    .D1(_1939_),
    .Y(_1940_));
 sky130_fd_sc_hd__nand4_2 _6167_ (.A(net299),
    .B(net224),
    .C(net218),
    .D(net307),
    .Y(_1941_));
 sky130_fd_sc_hd__a22o_1 _6168_ (.A1(net288),
    .A2(net229),
    .B1(_1939_),
    .B2(_1941_),
    .X(_1942_));
 sky130_fd_sc_hd__nand3b_4 _6169_ (.A_N(_1933_),
    .B(_1940_),
    .C(_1942_),
    .Y(_1943_));
 sky130_fd_sc_hd__o21ai_2 _6170_ (.A1(_1935_),
    .A2(_1936_),
    .B1(_1875_),
    .Y(_1944_));
 sky130_fd_sc_hd__o22a_2 _6171_ (.A1(_3022_),
    .A2(_1355_),
    .B1(_1415_),
    .B2(_2848_),
    .X(_1946_));
 sky130_fd_sc_hd__a21o_1 _6172_ (.A1(_1939_),
    .A2(_1941_),
    .B1(_1875_),
    .X(_1947_));
 sky130_fd_sc_hd__o211ai_4 _6173_ (.A1(_1944_),
    .A2(_1946_),
    .B1(_1933_),
    .C1(_1947_),
    .Y(_1948_));
 sky130_fd_sc_hd__a21boi_2 _6174_ (.A1(_1935_),
    .A2(_1823_),
    .B1_N(_1822_),
    .Y(_1949_));
 sky130_fd_sc_hd__a21oi_2 _6175_ (.A1(_1943_),
    .A2(_1948_),
    .B1(_1949_),
    .Y(_1950_));
 sky130_fd_sc_hd__and3_1 _6176_ (.A(_1949_),
    .B(_1943_),
    .C(_1948_),
    .X(_1951_));
 sky130_fd_sc_hd__inv_6 _6177_ (.A(net179),
    .Y(_1952_));
 sky130_fd_sc_hd__buf_6 _6178_ (.A(_1952_),
    .X(_1953_));
 sky130_fd_sc_hd__o2bb2ai_2 _6179_ (.A1_N(net370),
    .A2_N(net183),
    .B1(net389),
    .B2(_1953_),
    .Y(_1954_));
 sky130_fd_sc_hd__nand4_4 _6180_ (.A(_2982_),
    .B(net370),
    .C(net183),
    .D(net179),
    .Y(_1955_));
 sky130_fd_sc_hd__a21oi_4 _6181_ (.A1(_1954_),
    .A2(_1955_),
    .B1(_1848_),
    .Y(_1957_));
 sky130_fd_sc_hd__clkbuf_8 _6182_ (.A(_1952_),
    .X(_1958_));
 sky130_fd_sc_hd__a21oi_4 _6183_ (.A1(net388),
    .A2(net187),
    .B1(_3124_),
    .Y(_1959_));
 sky130_fd_sc_hd__nand3_1 _6184_ (.A(_1848_),
    .B(_1954_),
    .C(_1955_),
    .Y(_1960_));
 sky130_fd_sc_hd__o21ai_4 _6185_ (.A1(_1958_),
    .A2(_1959_),
    .B1(_1960_),
    .Y(_1961_));
 sky130_fd_sc_hd__a22oi_4 _6186_ (.A1(net370),
    .A2(net182),
    .B1(_2982_),
    .B2(net179),
    .Y(_1962_));
 sky130_fd_sc_hd__and4b_1 _6187_ (.A_N(net378),
    .B(net370),
    .C(net183),
    .D(net179),
    .X(_1963_));
 sky130_fd_sc_hd__o22ai_2 _6188_ (.A1(_1727_),
    .A2(_1642_),
    .B1(_1962_),
    .B2(_1963_),
    .Y(_1964_));
 sky130_fd_sc_hd__a21oi_1 _6189_ (.A1(_1732_),
    .A2(net392),
    .B1(_1958_),
    .Y(_1965_));
 sky130_fd_sc_hd__nand4_2 _6190_ (.A(_1954_),
    .B(_1955_),
    .C(net357),
    .D(net191),
    .Y(_1966_));
 sky130_fd_sc_hd__nand3_4 _6191_ (.A(_1964_),
    .B(_1965_),
    .C(_1966_),
    .Y(_1968_));
 sky130_fd_sc_hd__o21ai_1 _6192_ (.A1(_1957_),
    .A2(_1961_),
    .B1(_1968_),
    .Y(_1969_));
 sky130_fd_sc_hd__nand4_2 _6193_ (.A(net345),
    .B(net330),
    .C(net206),
    .D(net200),
    .Y(_1970_));
 sky130_fd_sc_hd__nand2_1 _6194_ (.A(net345),
    .B(net196),
    .Y(_1971_));
 sky130_fd_sc_hd__nand2_2 _6195_ (.A(net330),
    .B(net206),
    .Y(_1972_));
 sky130_fd_sc_hd__nand2_1 _6196_ (.A(net211),
    .B(net319),
    .Y(_1973_));
 sky130_fd_sc_hd__a21oi_1 _6197_ (.A1(_1971_),
    .A2(_1972_),
    .B1(_1973_),
    .Y(_1974_));
 sky130_fd_sc_hd__nand2_1 _6198_ (.A(_1971_),
    .B(_1972_),
    .Y(_1975_));
 sky130_fd_sc_hd__a22oi_2 _6199_ (.A1(net211),
    .A2(net318),
    .B1(_1975_),
    .B2(_1970_),
    .Y(_1976_));
 sky130_fd_sc_hd__a21oi_1 _6200_ (.A1(_1970_),
    .A2(_1974_),
    .B1(_1976_),
    .Y(_1977_));
 sky130_fd_sc_hd__nand2_1 _6201_ (.A(_1969_),
    .B(_1977_),
    .Y(_1979_));
 sky130_fd_sc_hd__o31a_1 _6202_ (.A1(net178),
    .A2(_1630_),
    .A3(_1732_),
    .B1(_1850_),
    .X(_1980_));
 sky130_fd_sc_hd__a21o_2 _6203_ (.A1(_1970_),
    .A2(_1974_),
    .B1(_1976_),
    .X(_1981_));
 sky130_fd_sc_hd__o211ai_2 _6204_ (.A1(_1957_),
    .A2(_1961_),
    .B1(_1981_),
    .C1(_1968_),
    .Y(_1982_));
 sky130_fd_sc_hd__nand3_4 _6205_ (.A(_1979_),
    .B(_1980_),
    .C(_1982_),
    .Y(_1983_));
 sky130_fd_sc_hd__inv_2 _6206_ (.A(_1850_),
    .Y(_1984_));
 sky130_fd_sc_hd__buf_6 _6207_ (.A(_1953_),
    .X(_1985_));
 sky130_fd_sc_hd__and4_1 _6208_ (.A(_1985_),
    .B(_1647_),
    .C(net378),
    .D(net183),
    .X(_1986_));
 sky130_fd_sc_hd__o211ai_2 _6209_ (.A1(_1957_),
    .A2(_1961_),
    .B1(_1977_),
    .C1(_1968_),
    .Y(_1987_));
 sky130_fd_sc_hd__nand2_1 _6210_ (.A(_1969_),
    .B(_1981_),
    .Y(_1988_));
 sky130_fd_sc_hd__o211ai_4 _6211_ (.A1(_1984_),
    .A2(_1986_),
    .B1(_1987_),
    .C1(_1988_),
    .Y(_1990_));
 sky130_fd_sc_hd__o211ai_2 _6212_ (.A1(_1950_),
    .A2(_1951_),
    .B1(_1983_),
    .C1(_1990_),
    .Y(_1991_));
 sky130_fd_sc_hd__a21boi_2 _6213_ (.A1(_1943_),
    .A2(_1948_),
    .B1_N(_1949_),
    .Y(_1992_));
 sky130_fd_sc_hd__and3b_1 _6214_ (.A_N(_1949_),
    .B(_1943_),
    .C(_1948_),
    .X(_1993_));
 sky130_fd_sc_hd__o2bb2ai_1 _6215_ (.A1_N(_1983_),
    .A2_N(_1990_),
    .B1(_1992_),
    .B2(_1993_),
    .Y(_1994_));
 sky130_fd_sc_hd__o211ai_4 _6216_ (.A1(_1928_),
    .A2(_1931_),
    .B1(_1991_),
    .C1(_1994_),
    .Y(_1995_));
 sky130_fd_sc_hd__o2bb2ai_1 _6217_ (.A1_N(_1983_),
    .A2_N(_1990_),
    .B1(_1950_),
    .B2(_1951_),
    .Y(_1996_));
 sky130_fd_sc_hd__o21ai_1 _6218_ (.A1(_1838_),
    .A2(_1928_),
    .B1(_1856_),
    .Y(_1997_));
 sky130_fd_sc_hd__o211ai_2 _6219_ (.A1(_1992_),
    .A2(_1993_),
    .B1(_1983_),
    .C1(_1990_),
    .Y(_1998_));
 sky130_fd_sc_hd__nand3_4 _6220_ (.A(_1996_),
    .B(_1997_),
    .C(_1998_),
    .Y(_1999_));
 sky130_fd_sc_hd__nor2_1 _6221_ (.A(_1835_),
    .B(_1832_),
    .Y(_2001_));
 sky130_fd_sc_hd__a22oi_1 _6222_ (.A1(net288),
    .A2(net234),
    .B1(net227),
    .B2(net300),
    .Y(_2002_));
 sky130_fd_sc_hd__o22ai_2 _6223_ (.A1(_1666_),
    .A2(_1875_),
    .B1(_1877_),
    .B2(_2002_),
    .Y(_2003_));
 sky130_fd_sc_hd__nand2_1 _6224_ (.A(net261),
    .B(net243),
    .Y(_2004_));
 sky130_fd_sc_hd__nand3_1 _6225_ (.A(_2004_),
    .B(net234),
    .C(net275),
    .Y(_2005_));
 sky130_fd_sc_hd__nand2_1 _6226_ (.A(net275),
    .B(net234),
    .Y(_2006_));
 sky130_fd_sc_hd__nand3_1 _6227_ (.A(_2006_),
    .B(net243),
    .C(net261),
    .Y(_2007_));
 sky130_fd_sc_hd__a21o_1 _6228_ (.A1(_2005_),
    .A2(_2007_),
    .B1(_1889_),
    .X(_2008_));
 sky130_fd_sc_hd__and2_1 _6229_ (.A(_2003_),
    .B(_2008_),
    .X(_2009_));
 sky130_fd_sc_hd__a22o_1 _6230_ (.A1(net261),
    .A2(net241),
    .B1(net234),
    .B2(net275),
    .X(_2010_));
 sky130_fd_sc_hd__nand4_1 _6231_ (.A(net275),
    .B(net261),
    .C(net241),
    .D(net234),
    .Y(_2012_));
 sky130_fd_sc_hd__nor2_4 _6232_ (.A(_1423_),
    .B(_1129_),
    .Y(_2013_));
 sky130_fd_sc_hd__a21o_1 _6233_ (.A1(_2010_),
    .A2(_2012_),
    .B1(_2013_),
    .X(_2014_));
 sky130_fd_sc_hd__a21oi_2 _6234_ (.A1(_2014_),
    .A2(_2008_),
    .B1(_2003_),
    .Y(_2015_));
 sky130_fd_sc_hd__a21oi_1 _6235_ (.A1(_2009_),
    .A2(_2014_),
    .B1(_2015_),
    .Y(_2016_));
 sky130_fd_sc_hd__o21ai_4 _6236_ (.A1(_1830_),
    .A2(_2001_),
    .B1(_2016_),
    .Y(_2017_));
 sky130_fd_sc_hd__and3_2 _6237_ (.A(_2008_),
    .B(_2003_),
    .C(_2014_),
    .X(_2018_));
 sky130_fd_sc_hd__o211ai_4 _6238_ (.A1(_2018_),
    .A2(_2015_),
    .B1(_1929_),
    .C1(_1930_),
    .Y(_2019_));
 sky130_fd_sc_hd__a21boi_4 _6239_ (.A1(_1883_),
    .A2(_2013_),
    .B1_N(_1887_),
    .Y(_2020_));
 sky130_fd_sc_hd__a21oi_2 _6240_ (.A1(_2017_),
    .A2(_2019_),
    .B1(_2020_),
    .Y(_2021_));
 sky130_fd_sc_hd__and3_1 _6241_ (.A(_2020_),
    .B(_2017_),
    .C(_2019_),
    .X(_2023_));
 sky130_fd_sc_hd__o2bb2ai_1 _6242_ (.A1_N(_1995_),
    .A2_N(_1999_),
    .B1(_2021_),
    .B2(_2023_),
    .Y(_2024_));
 sky130_fd_sc_hd__and3_2 _6243_ (.A(_1861_),
    .B(_1863_),
    .C(_1864_),
    .X(_2025_));
 sky130_fd_sc_hd__a31oi_2 _6244_ (.A1(_1870_),
    .A2(_1905_),
    .A3(_1899_),
    .B1(_2025_),
    .Y(_2026_));
 sky130_fd_sc_hd__and3b_1 _6245_ (.A_N(_2020_),
    .B(_2017_),
    .C(_2019_),
    .X(_2027_));
 sky130_fd_sc_hd__a21boi_2 _6246_ (.A1(_2017_),
    .A2(_2019_),
    .B1_N(_2020_),
    .Y(_2028_));
 sky130_fd_sc_hd__o211ai_2 _6247_ (.A1(_2027_),
    .A2(_2028_),
    .B1(_1995_),
    .C1(_1999_),
    .Y(_2029_));
 sky130_fd_sc_hd__nand3_1 _6248_ (.A(_2024_),
    .B(_2026_),
    .C(_2029_),
    .Y(_2030_));
 sky130_fd_sc_hd__o2111a_1 _6249_ (.A1(_1903_),
    .A2(_1904_),
    .B1(_1905_),
    .C1(_1865_),
    .D1(_1870_),
    .X(_2031_));
 sky130_fd_sc_hd__o211ai_2 _6250_ (.A1(_2021_),
    .A2(_2023_),
    .B1(_1995_),
    .C1(_1999_),
    .Y(_2032_));
 sky130_fd_sc_hd__o2bb2ai_1 _6251_ (.A1_N(_1995_),
    .A2_N(_1999_),
    .B1(_2027_),
    .B2(_2028_),
    .Y(_2034_));
 sky130_fd_sc_hd__o211ai_2 _6252_ (.A1(_2025_),
    .A2(_2031_),
    .B1(_2032_),
    .C1(_2034_),
    .Y(_2035_));
 sky130_fd_sc_hd__nand2_1 _6253_ (.A(_2030_),
    .B(_2035_),
    .Y(_2036_));
 sky130_fd_sc_hd__a32o_1 _6254_ (.A1(_1895_),
    .A2(_1893_),
    .A3(_1894_),
    .B1(_1892_),
    .B2(_1897_),
    .X(_2037_));
 sky130_fd_sc_hd__inv_2 _6255_ (.A(_2037_),
    .Y(_2038_));
 sky130_fd_sc_hd__nand2_1 _6256_ (.A(_2036_),
    .B(_2038_),
    .Y(_2039_));
 sky130_fd_sc_hd__nand3_1 _6257_ (.A(_2030_),
    .B(_2035_),
    .C(_2037_),
    .Y(_2040_));
 sky130_fd_sc_hd__nand2_1 _6258_ (.A(_2039_),
    .B(_2040_),
    .Y(_2041_));
 sky130_fd_sc_hd__o31a_2 _6259_ (.A1(_1715_),
    .A2(_1916_),
    .A3(_1917_),
    .B1(_1912_),
    .X(_2042_));
 sky130_fd_sc_hd__nand2_1 _6260_ (.A(_2041_),
    .B(_2042_),
    .Y(_2043_));
 sky130_fd_sc_hd__or2_1 _6261_ (.A(_2042_),
    .B(_2041_),
    .X(_2045_));
 sky130_fd_sc_hd__nand2_1 _6262_ (.A(_2043_),
    .B(_2045_),
    .Y(_2046_));
 sky130_fd_sc_hd__a32oi_4 _6263_ (.A1(_1919_),
    .A2(_1921_),
    .A3(_1915_),
    .B1(_1809_),
    .B2(_1810_),
    .Y(_2047_));
 sky130_fd_sc_hd__o211ai_4 _6264_ (.A1(_1606_),
    .A2(_1814_),
    .B1(_2047_),
    .C1(_1819_),
    .Y(_2048_));
 sky130_fd_sc_hd__o21bai_2 _6265_ (.A1(_1812_),
    .A2(_1922_),
    .B1_N(_1923_),
    .Y(_2049_));
 sky130_fd_sc_hd__nand2_2 _6266_ (.A(_2048_),
    .B(_2049_),
    .Y(_2050_));
 sky130_fd_sc_hd__xor2_1 _6267_ (.A(_2046_),
    .B(_2050_),
    .X(_0089_));
 sky130_fd_sc_hd__o211a_1 _6268_ (.A1(_2025_),
    .A2(_2031_),
    .B1(_2032_),
    .C1(_2034_),
    .X(_2051_));
 sky130_fd_sc_hd__a31oi_1 _6269_ (.A1(_2024_),
    .A2(_2026_),
    .A3(_2029_),
    .B1(_2038_),
    .Y(_2052_));
 sky130_fd_sc_hd__o21ai_1 _6270_ (.A1(_2027_),
    .A2(_2028_),
    .B1(_1999_),
    .Y(_2053_));
 sky130_fd_sc_hd__nand2_1 _6271_ (.A(_1995_),
    .B(_2053_),
    .Y(_2055_));
 sky130_fd_sc_hd__nand4_2 _6272_ (.A(net301),
    .B(net289),
    .C(net223),
    .D(net217),
    .Y(_2056_));
 sky130_fd_sc_hd__nand2_1 _6273_ (.A(net289),
    .B(net223),
    .Y(_2057_));
 sky130_fd_sc_hd__nand2_1 _6274_ (.A(_1936_),
    .B(_2057_),
    .Y(_2058_));
 sky130_fd_sc_hd__a22o_1 _6275_ (.A1(net276),
    .A2(net229),
    .B1(_2056_),
    .B2(_2058_),
    .X(_2059_));
 sky130_fd_sc_hd__nand2_1 _6276_ (.A(net289),
    .B(net218),
    .Y(_2060_));
 sky130_fd_sc_hd__o2111ai_1 _6277_ (.A1(_1938_),
    .A2(_2060_),
    .B1(net276),
    .C1(net229),
    .D1(_2058_),
    .Y(_2061_));
 sky130_fd_sc_hd__a22oi_2 _6278_ (.A1(_1971_),
    .A2(_1972_),
    .B1(_1970_),
    .B2(_1973_),
    .Y(_2062_));
 sky130_fd_sc_hd__nand3_2 _6279_ (.A(_2059_),
    .B(_2061_),
    .C(_2062_),
    .Y(_2063_));
 sky130_fd_sc_hd__o221ai_1 _6280_ (.A1(_2928_),
    .A2(_1331_),
    .B1(_1938_),
    .B2(_2060_),
    .C1(_2058_),
    .Y(_2064_));
 sky130_fd_sc_hd__o2bb2ai_1 _6281_ (.A1_N(_1936_),
    .A2_N(_2057_),
    .B1(_2060_),
    .B2(_1938_),
    .Y(_2066_));
 sky130_fd_sc_hd__nand3_1 _6282_ (.A(_2066_),
    .B(net229),
    .C(net277),
    .Y(_2067_));
 sky130_fd_sc_hd__nand3b_1 _6283_ (.A_N(_2062_),
    .B(_2064_),
    .C(_2067_),
    .Y(_2068_));
 sky130_fd_sc_hd__o21ai_1 _6284_ (.A1(_1875_),
    .A2(_1946_),
    .B1(_1941_),
    .Y(_2069_));
 sky130_fd_sc_hd__a21oi_1 _6285_ (.A1(_2063_),
    .A2(_2068_),
    .B1(_2069_),
    .Y(_2070_));
 sky130_fd_sc_hd__and3_1 _6286_ (.A(_2063_),
    .B(_2068_),
    .C(_2069_),
    .X(_2071_));
 sky130_fd_sc_hd__o21a_1 _6287_ (.A1(_1848_),
    .A2(_1962_),
    .B1(_1955_),
    .X(_2072_));
 sky130_fd_sc_hd__a22o_1 _6288_ (.A1(net353),
    .A2(net182),
    .B1(_2218_),
    .B2(net178),
    .X(_2073_));
 sky130_fd_sc_hd__nand4b_4 _6289_ (.A_N(net366),
    .B(net353),
    .C(net182),
    .D(net178),
    .Y(_2074_));
 sky130_fd_sc_hd__o211ai_2 _6290_ (.A1(_2965_),
    .A2(_1642_),
    .B1(_2073_),
    .C1(_2074_),
    .Y(_2075_));
 sky130_fd_sc_hd__a22oi_4 _6291_ (.A1(net354),
    .A2(net182),
    .B1(_2218_),
    .B2(net178),
    .Y(_2077_));
 sky130_fd_sc_hd__and4b_1 _6292_ (.A_N(net366),
    .B(net353),
    .C(net182),
    .D(net178),
    .X(_2078_));
 sky130_fd_sc_hd__nand2_2 _6293_ (.A(net341),
    .B(net191),
    .Y(_2079_));
 sky130_fd_sc_hd__o21bai_2 _6294_ (.A1(_2077_),
    .A2(_2078_),
    .B1_N(_2079_),
    .Y(_2080_));
 sky130_fd_sc_hd__nand3_4 _6295_ (.A(_2072_),
    .B(_2075_),
    .C(_2080_),
    .Y(_2081_));
 sky130_fd_sc_hd__o21ai_4 _6296_ (.A1(_2077_),
    .A2(_2078_),
    .B1(_2079_),
    .Y(_2082_));
 sky130_fd_sc_hd__nand4_4 _6297_ (.A(_2073_),
    .B(_2074_),
    .C(net341),
    .D(net191),
    .Y(_2083_));
 sky130_fd_sc_hd__o21ai_2 _6298_ (.A1(_1848_),
    .A2(_1962_),
    .B1(_1955_),
    .Y(_2084_));
 sky130_fd_sc_hd__nand3_4 _6299_ (.A(_2082_),
    .B(_2083_),
    .C(_2084_),
    .Y(_2085_));
 sky130_fd_sc_hd__nand2_1 _6300_ (.A(_2081_),
    .B(_2085_),
    .Y(_2086_));
 sky130_fd_sc_hd__a22oi_4 _6301_ (.A1(net319),
    .A2(net206),
    .B1(net196),
    .B2(net330),
    .Y(_2088_));
 sky130_fd_sc_hd__nand2_1 _6302_ (.A(net318),
    .B(net196),
    .Y(_2089_));
 sky130_fd_sc_hd__nor2_1 _6303_ (.A(_1972_),
    .B(_2089_),
    .Y(_2090_));
 sky130_fd_sc_hd__a21o_1 _6304_ (.A1(net211),
    .A2(net307),
    .B1(_2090_),
    .X(_2091_));
 sky130_fd_sc_hd__o211ai_2 _6305_ (.A1(_2088_),
    .A2(_2090_),
    .B1(net211),
    .C1(net307),
    .Y(_2092_));
 sky130_fd_sc_hd__o21ai_4 _6306_ (.A1(_2088_),
    .A2(_2091_),
    .B1(_2092_),
    .Y(_2093_));
 sky130_fd_sc_hd__nand2_2 _6307_ (.A(_2086_),
    .B(_2093_),
    .Y(_2094_));
 sky130_fd_sc_hd__o22a_1 _6308_ (.A1(_1394_),
    .A2(_2973_),
    .B1(_2088_),
    .B2(_2090_),
    .X(_2095_));
 sky130_fd_sc_hd__a22o_1 _6309_ (.A1(net318),
    .A2(net206),
    .B1(net196),
    .B2(net330),
    .X(_2096_));
 sky130_fd_sc_hd__o2111a_1 _6310_ (.A1(_1972_),
    .A2(_2089_),
    .B1(net210),
    .C1(net307),
    .D1(_2096_),
    .X(_2097_));
 sky130_fd_sc_hd__o211ai_4 _6311_ (.A1(_2095_),
    .A2(_2097_),
    .B1(_2081_),
    .C1(_2085_),
    .Y(_2099_));
 sky130_fd_sc_hd__o2bb2ai_4 _6312_ (.A1_N(_1981_),
    .A2_N(_1968_),
    .B1(_1957_),
    .B2(_1961_),
    .Y(_2100_));
 sky130_fd_sc_hd__nand3_2 _6313_ (.A(_2094_),
    .B(_2099_),
    .C(_2100_),
    .Y(_2101_));
 sky130_fd_sc_hd__a2bb2oi_2 _6314_ (.A1_N(_1957_),
    .A2_N(_1961_),
    .B1(_1981_),
    .B2(_1968_),
    .Y(_2102_));
 sky130_fd_sc_hd__nand3_1 _6315_ (.A(_2081_),
    .B(_2085_),
    .C(_2093_),
    .Y(_2103_));
 sky130_fd_sc_hd__o2bb2ai_2 _6316_ (.A1_N(_2081_),
    .A2_N(_2085_),
    .B1(_2095_),
    .B2(_2097_),
    .Y(_2104_));
 sky130_fd_sc_hd__nand3_1 _6317_ (.A(_2102_),
    .B(_2103_),
    .C(_2104_),
    .Y(_2105_));
 sky130_fd_sc_hd__o211ai_1 _6318_ (.A1(_2070_),
    .A2(_2071_),
    .B1(_2101_),
    .C1(_2105_),
    .Y(_2106_));
 sky130_fd_sc_hd__nand2_1 _6319_ (.A(_2105_),
    .B(_2101_),
    .Y(_2107_));
 sky130_fd_sc_hd__nor2_1 _6320_ (.A(_2070_),
    .B(_2071_),
    .Y(_2108_));
 sky130_fd_sc_hd__nand2_1 _6321_ (.A(_2107_),
    .B(_2108_),
    .Y(_2110_));
 sky130_fd_sc_hd__o21ai_1 _6322_ (.A1(_1950_),
    .A2(_1951_),
    .B1(_1990_),
    .Y(_2111_));
 sky130_fd_sc_hd__nand2_2 _6323_ (.A(_1983_),
    .B(_2111_),
    .Y(_2112_));
 sky130_fd_sc_hd__nand3_2 _6324_ (.A(_2106_),
    .B(_2110_),
    .C(_2112_),
    .Y(_2113_));
 sky130_fd_sc_hd__nand2_1 _6325_ (.A(_2101_),
    .B(_2108_),
    .Y(_2114_));
 sky130_fd_sc_hd__a21oi_2 _6326_ (.A1(_2094_),
    .A2(_2099_),
    .B1(_2100_),
    .Y(_2115_));
 sky130_fd_sc_hd__nor2_1 _6327_ (.A(_1992_),
    .B(_1993_),
    .Y(_2116_));
 sky130_fd_sc_hd__a21boi_2 _6328_ (.A1(_1990_),
    .A2(_2116_),
    .B1_N(_1983_),
    .Y(_2117_));
 sky130_fd_sc_hd__a21o_1 _6329_ (.A1(_2105_),
    .A2(_2101_),
    .B1(_2108_),
    .X(_2118_));
 sky130_fd_sc_hd__o211ai_2 _6330_ (.A1(_2114_),
    .A2(_2115_),
    .B1(_2117_),
    .C1(_2118_),
    .Y(_2119_));
 sky130_fd_sc_hd__nand2_1 _6331_ (.A(_1949_),
    .B(_1948_),
    .Y(_2121_));
 sky130_fd_sc_hd__nand3_1 _6332_ (.A(net261),
    .B(net241),
    .C(net236),
    .Y(_2122_));
 sky130_fd_sc_hd__o21a_1 _6333_ (.A1(net241),
    .A2(net235),
    .B1(net265),
    .X(_2123_));
 sky130_fd_sc_hd__buf_2 _6334_ (.A(_2123_),
    .X(_2124_));
 sky130_fd_sc_hd__o211ai_1 _6335_ (.A1(_1889_),
    .A2(_2010_),
    .B1(_2122_),
    .C1(_2124_),
    .Y(_2125_));
 sky130_fd_sc_hd__a211o_1 _6336_ (.A1(_2123_),
    .A2(_2122_),
    .B1(_1301_),
    .C1(_3058_),
    .X(_2126_));
 sky130_fd_sc_hd__and4_1 _6337_ (.A(net265),
    .B(net249),
    .C(net241),
    .D(net235),
    .X(_2127_));
 sky130_fd_sc_hd__a31o_1 _6338_ (.A1(_2012_),
    .A2(_2125_),
    .A3(_2126_),
    .B1(_2127_),
    .X(_2128_));
 sky130_fd_sc_hd__nand3_1 _6339_ (.A(_1943_),
    .B(_2121_),
    .C(_2128_),
    .Y(_2129_));
 sky130_fd_sc_hd__a21o_1 _6340_ (.A1(_1943_),
    .A2(_2121_),
    .B1(_2128_),
    .X(_2130_));
 sky130_fd_sc_hd__nand2_1 _6341_ (.A(_2009_),
    .B(_2014_),
    .Y(_2132_));
 sky130_fd_sc_hd__a21oi_1 _6342_ (.A1(_2129_),
    .A2(_2130_),
    .B1(_2132_),
    .Y(_2133_));
 sky130_fd_sc_hd__and3_1 _6343_ (.A(_2132_),
    .B(_2129_),
    .C(_2130_),
    .X(_2134_));
 sky130_fd_sc_hd__o2bb2ai_1 _6344_ (.A1_N(_2113_),
    .A2_N(_2119_),
    .B1(_2133_),
    .B2(_2134_),
    .Y(_2135_));
 sky130_fd_sc_hd__and3_1 _6345_ (.A(_2130_),
    .B(_2018_),
    .C(_2129_),
    .X(_2136_));
 sky130_fd_sc_hd__a21oi_1 _6346_ (.A1(_2129_),
    .A2(_2130_),
    .B1(_2018_),
    .Y(_2137_));
 sky130_fd_sc_hd__o211ai_1 _6347_ (.A1(_2136_),
    .A2(_2137_),
    .B1(_2113_),
    .C1(_2119_),
    .Y(_2138_));
 sky130_fd_sc_hd__nand3_2 _6348_ (.A(_2055_),
    .B(_2135_),
    .C(_2138_),
    .Y(_2139_));
 sky130_fd_sc_hd__o2bb2ai_1 _6349_ (.A1_N(_2113_),
    .A2_N(_2119_),
    .B1(_2136_),
    .B2(_2137_),
    .Y(_2140_));
 sky130_fd_sc_hd__o211ai_1 _6350_ (.A1(_2133_),
    .A2(_2134_),
    .B1(_2113_),
    .C1(_2119_),
    .Y(_2141_));
 sky130_fd_sc_hd__o21ai_1 _6351_ (.A1(_2021_),
    .A2(_2023_),
    .B1(_1995_),
    .Y(_2143_));
 sky130_fd_sc_hd__nand2_1 _6352_ (.A(_1999_),
    .B(_2143_),
    .Y(_2144_));
 sky130_fd_sc_hd__nand3_2 _6353_ (.A(_2140_),
    .B(_2141_),
    .C(_2144_),
    .Y(_2145_));
 sky130_fd_sc_hd__o211a_1 _6354_ (.A1(_2018_),
    .A2(_2015_),
    .B1(_1929_),
    .C1(_1834_),
    .X(_2146_));
 sky130_fd_sc_hd__o21ai_2 _6355_ (.A1(_2020_),
    .A2(_2146_),
    .B1(_2017_),
    .Y(_2147_));
 sky130_fd_sc_hd__nand3_1 _6356_ (.A(_2139_),
    .B(_2145_),
    .C(_2147_),
    .Y(_2148_));
 sky130_fd_sc_hd__a21o_1 _6357_ (.A1(_2139_),
    .A2(_2145_),
    .B1(_2147_),
    .X(_2149_));
 sky130_fd_sc_hd__o211ai_2 _6358_ (.A1(_2051_),
    .A2(_2052_),
    .B1(_2148_),
    .C1(_2149_),
    .Y(_2150_));
 sky130_fd_sc_hd__nand2_1 _6359_ (.A(_2139_),
    .B(_2145_),
    .Y(_2151_));
 sky130_fd_sc_hd__nand2_1 _6360_ (.A(_2151_),
    .B(_2147_),
    .Y(_2152_));
 sky130_fd_sc_hd__o21ai_1 _6361_ (.A1(_2037_),
    .A2(_2051_),
    .B1(_2030_),
    .Y(_2154_));
 sky130_fd_sc_hd__o2111ai_2 _6362_ (.A1(_2146_),
    .A2(_2020_),
    .B1(_2017_),
    .C1(_2139_),
    .D1(_2145_),
    .Y(_2155_));
 sky130_fd_sc_hd__nand3_2 _6363_ (.A(_2152_),
    .B(_2154_),
    .C(_2155_),
    .Y(_2156_));
 sky130_fd_sc_hd__o21ai_1 _6364_ (.A1(_2050_),
    .A2(_2046_),
    .B1(_2045_),
    .Y(_2157_));
 sky130_fd_sc_hd__a21oi_1 _6365_ (.A1(_2150_),
    .A2(_2156_),
    .B1(_2157_),
    .Y(_2158_));
 sky130_fd_sc_hd__and3_1 _6366_ (.A(_2150_),
    .B(_2156_),
    .C(_2157_),
    .X(_2159_));
 sky130_fd_sc_hd__nor2_1 _6367_ (.A(_2158_),
    .B(_2159_),
    .Y(_0090_));
 sky130_fd_sc_hd__o21ai_1 _6368_ (.A1(_2115_),
    .A2(_2114_),
    .B1(_2118_),
    .Y(_2160_));
 sky130_fd_sc_hd__o21ai_1 _6369_ (.A1(_2133_),
    .A2(_2134_),
    .B1(_2113_),
    .Y(_2161_));
 sky130_fd_sc_hd__o21ai_1 _6370_ (.A1(_2160_),
    .A2(_2112_),
    .B1(_2161_),
    .Y(_2162_));
 sky130_fd_sc_hd__a22o_1 _6371_ (.A1(_1939_),
    .A2(_1944_),
    .B1(_2063_),
    .B2(_2068_),
    .X(_2164_));
 sky130_fd_sc_hd__nand4_1 _6372_ (.A(_1939_),
    .B(_1944_),
    .C(_2063_),
    .D(_2068_),
    .Y(_2165_));
 sky130_fd_sc_hd__nand2_1 _6373_ (.A(_2164_),
    .B(_2165_),
    .Y(_2166_));
 sky130_fd_sc_hd__a31oi_2 _6374_ (.A1(_2100_),
    .A2(_2094_),
    .A3(_2099_),
    .B1(_2166_),
    .Y(_2167_));
 sky130_fd_sc_hd__a31o_1 _6375_ (.A1(_2096_),
    .A2(net307),
    .A3(net210),
    .B1(_2090_),
    .X(_2168_));
 sky130_fd_sc_hd__nand4_2 _6376_ (.A(net289),
    .B(net276),
    .C(net223),
    .D(net217),
    .Y(_2169_));
 sky130_fd_sc_hd__a22o_1 _6377_ (.A1(net276),
    .A2(net223),
    .B1(net217),
    .B2(net289),
    .X(_2170_));
 sky130_fd_sc_hd__a22o_1 _6378_ (.A1(net262),
    .A2(net229),
    .B1(_2169_),
    .B2(_2170_),
    .X(_2171_));
 sky130_fd_sc_hd__nand4_1 _6379_ (.A(_2170_),
    .B(net230),
    .C(net262),
    .D(_2169_),
    .Y(_2172_));
 sky130_fd_sc_hd__nand3_2 _6380_ (.A(_2168_),
    .B(_2171_),
    .C(_2172_),
    .Y(_2173_));
 sky130_fd_sc_hd__o22a_1 _6381_ (.A1(_1393_),
    .A2(_2973_),
    .B1(_1972_),
    .B2(_2089_),
    .X(_2175_));
 sky130_fd_sc_hd__o211ai_2 _6382_ (.A1(_3058_),
    .A2(_1331_),
    .B1(_2169_),
    .C1(_2170_),
    .Y(_2176_));
 sky130_fd_sc_hd__nand2_4 _6383_ (.A(net262),
    .B(net230),
    .Y(_2177_));
 sky130_fd_sc_hd__a21o_1 _6384_ (.A1(_2169_),
    .A2(_2170_),
    .B1(_2177_),
    .X(_2178_));
 sky130_fd_sc_hd__o211ai_4 _6385_ (.A1(_2088_),
    .A2(_2175_),
    .B1(_2176_),
    .C1(_2178_),
    .Y(_2179_));
 sky130_fd_sc_hd__nand2_1 _6386_ (.A(net277),
    .B(net229),
    .Y(_2180_));
 sky130_fd_sc_hd__a22o_1 _6387_ (.A1(_2180_),
    .A2(_2056_),
    .B1(_2057_),
    .B2(_1936_),
    .X(_2181_));
 sky130_fd_sc_hd__a21oi_1 _6388_ (.A1(_2173_),
    .A2(_2179_),
    .B1(_2181_),
    .Y(_2182_));
 sky130_fd_sc_hd__and3_1 _6389_ (.A(_2173_),
    .B(_2179_),
    .C(_2181_),
    .X(_2183_));
 sky130_fd_sc_hd__a22o_1 _6390_ (.A1(net206),
    .A2(net314),
    .B1(net196),
    .B2(net326),
    .X(_2184_));
 sky130_fd_sc_hd__nand4_1 _6391_ (.A(net318),
    .B(net206),
    .C(net307),
    .D(net196),
    .Y(_2186_));
 sky130_fd_sc_hd__a22o_1 _6392_ (.A1(net301),
    .A2(net210),
    .B1(_2184_),
    .B2(_2186_),
    .X(_2187_));
 sky130_fd_sc_hd__nand4_2 _6393_ (.A(_2184_),
    .B(_2186_),
    .C(net301),
    .D(net210),
    .Y(_2188_));
 sky130_fd_sc_hd__nand2_2 _6394_ (.A(_2187_),
    .B(_2188_),
    .Y(_2189_));
 sky130_fd_sc_hd__inv_2 _6395_ (.A(_2189_),
    .Y(_2190_));
 sky130_fd_sc_hd__o2bb2ai_1 _6396_ (.A1_N(net340),
    .A2_N(net184),
    .B1(net359),
    .B2(_1952_),
    .Y(_2191_));
 sky130_fd_sc_hd__buf_4 _6397_ (.A(_2191_),
    .X(_2192_));
 sky130_fd_sc_hd__nand4b_4 _6398_ (.A_N(net359),
    .B(net340),
    .C(net184),
    .D(net179),
    .Y(_2193_));
 sky130_fd_sc_hd__and2_2 _6399_ (.A(net332),
    .B(net191),
    .X(_2194_));
 sky130_fd_sc_hd__a21oi_1 _6400_ (.A1(_2192_),
    .A2(_2193_),
    .B1(_2194_),
    .Y(_2195_));
 sky130_fd_sc_hd__and2_1 _6401_ (.A(net357),
    .B(net184),
    .X(_2197_));
 sky130_fd_sc_hd__nor2_1 _6402_ (.A(net370),
    .B(_1985_),
    .Y(_2198_));
 sky130_fd_sc_hd__clkbuf_4 _6403_ (.A(_1641_),
    .X(_2199_));
 sky130_fd_sc_hd__o21ai_1 _6404_ (.A1(_0385_),
    .A2(_2199_),
    .B1(_2074_),
    .Y(_2200_));
 sky130_fd_sc_hd__nand3_2 _6405_ (.A(_2192_),
    .B(_2193_),
    .C(_2194_),
    .Y(_2201_));
 sky130_fd_sc_hd__o211ai_1 _6406_ (.A1(_2197_),
    .A2(_2198_),
    .B1(_2200_),
    .C1(_2201_),
    .Y(_2202_));
 sky130_fd_sc_hd__nand3_1 _6407_ (.A(_1727_),
    .B(net341),
    .C(net184),
    .Y(_2203_));
 sky130_fd_sc_hd__o221a_2 _6408_ (.A1(_3441_),
    .A2(_2199_),
    .B1(_1985_),
    .B2(_2203_),
    .C1(_2192_),
    .X(_2204_));
 sky130_fd_sc_hd__nand2_1 _6409_ (.A(_2192_),
    .B(_2193_),
    .Y(_2205_));
 sky130_fd_sc_hd__o21a_1 _6410_ (.A1(_2965_),
    .A2(_1642_),
    .B1(_2074_),
    .X(_2206_));
 sky130_fd_sc_hd__o2bb2ai_4 _6411_ (.A1_N(_2194_),
    .A2_N(_2205_),
    .B1(_2077_),
    .B2(_2206_),
    .Y(_2208_));
 sky130_fd_sc_hd__o22ai_1 _6412_ (.A1(_2195_),
    .A2(_2202_),
    .B1(_2204_),
    .B2(_2208_),
    .Y(_2209_));
 sky130_fd_sc_hd__nand2_1 _6413_ (.A(_2190_),
    .B(_2209_),
    .Y(_2210_));
 sky130_fd_sc_hd__a32oi_4 _6414_ (.A1(_2084_),
    .A2(_2082_),
    .A3(_2083_),
    .B1(_2081_),
    .B2(_2093_),
    .Y(_2211_));
 sky130_fd_sc_hd__a22o_1 _6415_ (.A1(net332),
    .A2(net190),
    .B1(_2192_),
    .B2(_2193_),
    .X(_2212_));
 sky130_fd_sc_hd__o21ai_2 _6416_ (.A1(_2079_),
    .A2(_2077_),
    .B1(_2074_),
    .Y(_2213_));
 sky130_fd_sc_hd__nand3_4 _6417_ (.A(_2212_),
    .B(_2201_),
    .C(_2213_),
    .Y(_2214_));
 sky130_fd_sc_hd__o211ai_2 _6418_ (.A1(_2204_),
    .A2(_2208_),
    .B1(_2189_),
    .C1(_2214_),
    .Y(_2215_));
 sky130_fd_sc_hd__nand3_4 _6419_ (.A(_2210_),
    .B(_2211_),
    .C(_2215_),
    .Y(_2216_));
 sky130_fd_sc_hd__nand2_1 _6420_ (.A(_2081_),
    .B(_2093_),
    .Y(_2217_));
 sky130_fd_sc_hd__nand2_1 _6421_ (.A(_2085_),
    .B(_2217_),
    .Y(_2219_));
 sky130_fd_sc_hd__o2111ai_4 _6422_ (.A1(_2204_),
    .A2(_2208_),
    .B1(_2187_),
    .C1(_2188_),
    .D1(_2214_),
    .Y(_2220_));
 sky130_fd_sc_hd__nand2_1 _6423_ (.A(_2209_),
    .B(_2189_),
    .Y(_2221_));
 sky130_fd_sc_hd__nand3_4 _6424_ (.A(_2219_),
    .B(_2220_),
    .C(_2221_),
    .Y(_2222_));
 sky130_fd_sc_hd__o211ai_2 _6425_ (.A1(_2182_),
    .A2(_2183_),
    .B1(_2216_),
    .C1(_2222_),
    .Y(_2223_));
 sky130_fd_sc_hd__a22oi_2 _6426_ (.A1(_2180_),
    .A2(_2056_),
    .B1(_2057_),
    .B2(_1936_),
    .Y(_2224_));
 sky130_fd_sc_hd__a21oi_2 _6427_ (.A1(_2173_),
    .A2(_2179_),
    .B1(_2224_),
    .Y(_2225_));
 sky130_fd_sc_hd__and3_1 _6428_ (.A(_2173_),
    .B(_2179_),
    .C(_2224_),
    .X(_2226_));
 sky130_fd_sc_hd__o2bb2ai_2 _6429_ (.A1_N(_2216_),
    .A2_N(_2222_),
    .B1(_2225_),
    .B2(_2226_),
    .Y(_2227_));
 sky130_fd_sc_hd__o211ai_4 _6430_ (.A1(_2115_),
    .A2(_2167_),
    .B1(_2223_),
    .C1(_2227_),
    .Y(_2228_));
 sky130_fd_sc_hd__o2bb2ai_1 _6431_ (.A1_N(_2216_),
    .A2_N(_2222_),
    .B1(_2182_),
    .B2(_2183_),
    .Y(_2230_));
 sky130_fd_sc_hd__a32oi_2 _6432_ (.A1(_2102_),
    .A2(_2103_),
    .A3(_2104_),
    .B1(_2101_),
    .B2(_2108_),
    .Y(_2231_));
 sky130_fd_sc_hd__o211ai_1 _6433_ (.A1(_2225_),
    .A2(_2226_),
    .B1(_2216_),
    .C1(_2222_),
    .Y(_2232_));
 sky130_fd_sc_hd__nand3_2 _6434_ (.A(_2230_),
    .B(_2231_),
    .C(_2232_),
    .Y(_2233_));
 sky130_fd_sc_hd__a21oi_2 _6435_ (.A1(net264),
    .A2(net251),
    .B1(_2124_),
    .Y(_2234_));
 sky130_fd_sc_hd__and3_1 _6436_ (.A(_2063_),
    .B(_2165_),
    .C(_2234_),
    .X(_2235_));
 sky130_fd_sc_hd__o2bb2a_2 _6437_ (.A1_N(_2063_),
    .A2_N(_2165_),
    .B1(_2124_),
    .B2(_2013_),
    .X(_2236_));
 sky130_fd_sc_hd__nor2_1 _6438_ (.A(_2235_),
    .B(_2236_),
    .Y(_2237_));
 sky130_fd_sc_hd__nand3_1 _6439_ (.A(_2228_),
    .B(_2233_),
    .C(_2237_),
    .Y(_2238_));
 sky130_fd_sc_hd__a21o_1 _6440_ (.A1(_2228_),
    .A2(_2233_),
    .B1(_2237_),
    .X(_2239_));
 sky130_fd_sc_hd__and3_1 _6441_ (.A(_2162_),
    .B(_2238_),
    .C(_2239_),
    .X(_2241_));
 sky130_fd_sc_hd__o211ai_1 _6442_ (.A1(_2235_),
    .A2(_2236_),
    .B1(_2228_),
    .C1(_2233_),
    .Y(_2242_));
 sky130_fd_sc_hd__nand2_1 _6443_ (.A(_2228_),
    .B(_2233_),
    .Y(_2243_));
 sky130_fd_sc_hd__nand2_1 _6444_ (.A(_2243_),
    .B(_2237_),
    .Y(_2244_));
 sky130_fd_sc_hd__o2111ai_2 _6445_ (.A1(_2160_),
    .A2(_2112_),
    .B1(_2161_),
    .C1(_2242_),
    .D1(_2244_),
    .Y(_2245_));
 sky130_fd_sc_hd__a21bo_1 _6446_ (.A1(_2018_),
    .A2(_2129_),
    .B1_N(_2130_),
    .X(_2246_));
 sky130_fd_sc_hd__nand2_1 _6447_ (.A(_2245_),
    .B(_2246_),
    .Y(_2247_));
 sky130_fd_sc_hd__nand3_1 _6448_ (.A(_2162_),
    .B(_2238_),
    .C(_2239_),
    .Y(_2248_));
 sky130_fd_sc_hd__a21o_1 _6449_ (.A1(_2248_),
    .A2(_2245_),
    .B1(_2246_),
    .X(_2249_));
 sky130_fd_sc_hd__o21ai_1 _6450_ (.A1(_2241_),
    .A2(_2247_),
    .B1(_2249_),
    .Y(_2250_));
 sky130_fd_sc_hd__a21boi_1 _6451_ (.A1(_2139_),
    .A2(_2147_),
    .B1_N(_2145_),
    .Y(_2252_));
 sky130_fd_sc_hd__nand2_1 _6452_ (.A(_2250_),
    .B(_2252_),
    .Y(_2253_));
 sky130_fd_sc_hd__a21bo_1 _6453_ (.A1(_2147_),
    .A2(_2139_),
    .B1_N(_2145_),
    .X(_2254_));
 sky130_fd_sc_hd__o211ai_2 _6454_ (.A1(_2241_),
    .A2(_2247_),
    .B1(_2249_),
    .C1(_2254_),
    .Y(_2255_));
 sky130_fd_sc_hd__nand2_1 _6455_ (.A(_2253_),
    .B(_2255_),
    .Y(_2256_));
 sky130_fd_sc_hd__o21ai_1 _6456_ (.A1(_2042_),
    .A2(_2041_),
    .B1(_2150_),
    .Y(_2257_));
 sky130_fd_sc_hd__o211a_1 _6457_ (.A1(_2042_),
    .A2(_2041_),
    .B1(_2156_),
    .C1(_2150_),
    .X(_2258_));
 sky130_fd_sc_hd__nand2_1 _6458_ (.A(_2258_),
    .B(_2043_),
    .Y(_2259_));
 sky130_fd_sc_hd__o2bb2ai_1 _6459_ (.A1_N(_2156_),
    .A2_N(_2257_),
    .B1(_2050_),
    .B2(_2259_),
    .Y(_2260_));
 sky130_fd_sc_hd__xnor2_1 _6460_ (.A(_2256_),
    .B(_2260_),
    .Y(_0091_));
 sky130_fd_sc_hd__a21boi_1 _6461_ (.A1(_2233_),
    .A2(_2237_),
    .B1_N(_2228_),
    .Y(_2262_));
 sky130_fd_sc_hd__a32o_1 _6462_ (.A1(_2168_),
    .A2(_2171_),
    .A3(_2172_),
    .B1(_2179_),
    .B2(_2224_),
    .X(_2263_));
 sky130_fd_sc_hd__o311a_1 _6463_ (.A1(net251),
    .A2(net244),
    .A3(net236),
    .B1(_2263_),
    .C1(net263),
    .X(_2264_));
 sky130_fd_sc_hd__a211oi_1 _6464_ (.A1(net263),
    .A2(net251),
    .B1(_2124_),
    .C1(_2263_),
    .Y(_2265_));
 sky130_fd_sc_hd__o21ai_1 _6465_ (.A1(_2120_),
    .A2(_1642_),
    .B1(_2193_),
    .Y(_2266_));
 sky130_fd_sc_hd__nand2_1 _6466_ (.A(_2192_),
    .B(_2266_),
    .Y(_2267_));
 sky130_fd_sc_hd__o2bb2ai_2 _6467_ (.A1_N(net333),
    .A2_N(net185),
    .B1(net347),
    .B2(_1953_),
    .Y(_2268_));
 sky130_fd_sc_hd__nand4_4 _6468_ (.A(_1825_),
    .B(net333),
    .C(net185),
    .D(net180),
    .Y(_2269_));
 sky130_fd_sc_hd__o211ai_4 _6469_ (.A1(_2886_),
    .A2(_2199_),
    .B1(_2268_),
    .C1(_2269_),
    .Y(_2270_));
 sky130_fd_sc_hd__a22oi_4 _6470_ (.A1(net338),
    .A2(net186),
    .B1(_2965_),
    .B2(net179),
    .Y(_2271_));
 sky130_fd_sc_hd__and4b_1 _6471_ (.A_N(net351),
    .B(net338),
    .C(net184),
    .D(net181),
    .X(_2273_));
 sky130_fd_sc_hd__nor2_1 _6472_ (.A(_2886_),
    .B(_1642_),
    .Y(_2274_));
 sky130_fd_sc_hd__o21ai_2 _6473_ (.A1(_2271_),
    .A2(_2273_),
    .B1(_2274_),
    .Y(_2275_));
 sky130_fd_sc_hd__nand3_2 _6474_ (.A(_2267_),
    .B(_2270_),
    .C(_2275_),
    .Y(_2276_));
 sky130_fd_sc_hd__nand2_2 _6475_ (.A(net326),
    .B(net192),
    .Y(_2277_));
 sky130_fd_sc_hd__o21ai_2 _6476_ (.A1(_2271_),
    .A2(_2273_),
    .B1(_2277_),
    .Y(_2278_));
 sky130_fd_sc_hd__nand4_2 _6477_ (.A(_2268_),
    .B(_2269_),
    .C(net324),
    .D(net194),
    .Y(_2279_));
 sky130_fd_sc_hd__o2bb2ai_2 _6478_ (.A1_N(_2194_),
    .A2_N(_2191_),
    .B1(_2203_),
    .B2(_1958_),
    .Y(_2280_));
 sky130_fd_sc_hd__nand3_4 _6479_ (.A(_2278_),
    .B(_2279_),
    .C(_2280_),
    .Y(_2281_));
 sky130_fd_sc_hd__nand4_1 _6480_ (.A(net303),
    .B(net204),
    .C(net313),
    .D(net198),
    .Y(_2282_));
 sky130_fd_sc_hd__clkbuf_2 _6481_ (.A(_2282_),
    .X(_2284_));
 sky130_fd_sc_hd__a22o_2 _6482_ (.A1(net303),
    .A2(net206),
    .B1(net313),
    .B2(net196),
    .X(_2285_));
 sky130_fd_sc_hd__a22oi_2 _6483_ (.A1(net293),
    .A2(net210),
    .B1(_2284_),
    .B2(_2285_),
    .Y(_2286_));
 sky130_fd_sc_hd__and4_1 _6484_ (.A(_2285_),
    .B(net210),
    .C(net293),
    .D(_2284_),
    .X(_2287_));
 sky130_fd_sc_hd__nor2_1 _6485_ (.A(_2286_),
    .B(_2287_),
    .Y(_2288_));
 sky130_fd_sc_hd__a21o_1 _6486_ (.A1(_2276_),
    .A2(_2281_),
    .B1(_2288_),
    .X(_2289_));
 sky130_fd_sc_hd__a2bb2oi_2 _6487_ (.A1_N(_2204_),
    .A2_N(_2208_),
    .B1(_2189_),
    .B2(_2214_),
    .Y(_2290_));
 sky130_fd_sc_hd__a22o_1 _6488_ (.A1(net290),
    .A2(net213),
    .B1(_2284_),
    .B2(_2285_),
    .X(_2291_));
 sky130_fd_sc_hd__nand4_2 _6489_ (.A(_2285_),
    .B(net213),
    .C(net290),
    .D(_2284_),
    .Y(_2292_));
 sky130_fd_sc_hd__nand4_2 _6490_ (.A(_2276_),
    .B(_2281_),
    .C(_2291_),
    .D(_2292_),
    .Y(_2293_));
 sky130_fd_sc_hd__nand3_4 _6491_ (.A(_2289_),
    .B(_2290_),
    .C(_2293_),
    .Y(_2295_));
 sky130_fd_sc_hd__o21ai_2 _6492_ (.A1(_2286_),
    .A2(_2287_),
    .B1(_2281_),
    .Y(_2296_));
 sky130_fd_sc_hd__and3_1 _6493_ (.A(_2267_),
    .B(_2270_),
    .C(_2275_),
    .X(_2297_));
 sky130_fd_sc_hd__o2bb2ai_1 _6494_ (.A1_N(_2189_),
    .A2_N(_2214_),
    .B1(_2204_),
    .B2(_2208_),
    .Y(_2298_));
 sky130_fd_sc_hd__nand2_1 _6495_ (.A(net290),
    .B(net212),
    .Y(_2299_));
 sky130_fd_sc_hd__and3_1 _6496_ (.A(_2299_),
    .B(_2284_),
    .C(_2285_),
    .X(_2300_));
 sky130_fd_sc_hd__a21oi_1 _6497_ (.A1(_2284_),
    .A2(_2285_),
    .B1(_2299_),
    .Y(_2301_));
 sky130_fd_sc_hd__o2bb2ai_2 _6498_ (.A1_N(_2276_),
    .A2_N(_2281_),
    .B1(_2300_),
    .B2(_2301_),
    .Y(_2302_));
 sky130_fd_sc_hd__o211ai_4 _6499_ (.A1(_2296_),
    .A2(_2297_),
    .B1(_2298_),
    .C1(_2302_),
    .Y(_2303_));
 sky130_fd_sc_hd__nand4_4 _6500_ (.A(net276),
    .B(net262),
    .C(net222),
    .D(net216),
    .Y(_2304_));
 sky130_fd_sc_hd__o21ai_1 _6501_ (.A1(_3342_),
    .A2(_1331_),
    .B1(_2304_),
    .Y(_2306_));
 sky130_fd_sc_hd__o22a_2 _6502_ (.A1(_1423_),
    .A2(_1355_),
    .B1(_1415_),
    .B2(_2928_),
    .X(_2307_));
 sky130_fd_sc_hd__and4_1 _6503_ (.A(net326),
    .B(net206),
    .C(net314),
    .D(net196),
    .X(_2308_));
 sky130_fd_sc_hd__a31oi_1 _6504_ (.A1(_2184_),
    .A2(net210),
    .A3(net303),
    .B1(_2308_),
    .Y(_2309_));
 sky130_fd_sc_hd__a22o_1 _6505_ (.A1(net262),
    .A2(net222),
    .B1(net217),
    .B2(net276),
    .X(_2310_));
 sky130_fd_sc_hd__a21o_1 _6506_ (.A1(_2310_),
    .A2(_2304_),
    .B1(_2177_),
    .X(_2311_));
 sky130_fd_sc_hd__o211ai_2 _6507_ (.A1(_2306_),
    .A2(_2307_),
    .B1(_2309_),
    .C1(_2311_),
    .Y(_2312_));
 sky130_fd_sc_hd__and4_1 _6508_ (.A(net289),
    .B(net276),
    .C(net222),
    .D(net216),
    .X(_2313_));
 sky130_fd_sc_hd__a31o_1 _6509_ (.A1(_2170_),
    .A2(net230),
    .A3(net262),
    .B1(_2313_),
    .X(_2314_));
 sky130_fd_sc_hd__and2_1 _6510_ (.A(_2312_),
    .B(_2314_),
    .X(_2315_));
 sky130_fd_sc_hd__a41o_1 _6511_ (.A1(net276),
    .A2(net262),
    .A3(net222),
    .A4(net216),
    .B1(_2177_),
    .X(_2317_));
 sky130_fd_sc_hd__a22o_1 _6512_ (.A1(net262),
    .A2(net230),
    .B1(_2310_),
    .B2(_2304_),
    .X(_2318_));
 sky130_fd_sc_hd__a31o_1 _6513_ (.A1(_2184_),
    .A2(net210),
    .A3(net304),
    .B1(_2308_),
    .X(_2319_));
 sky130_fd_sc_hd__o211ai_4 _6514_ (.A1(_2307_),
    .A2(_2317_),
    .B1(_2318_),
    .C1(_2319_),
    .Y(_2320_));
 sky130_fd_sc_hd__a21oi_1 _6515_ (.A1(_2312_),
    .A2(_2320_),
    .B1(_2314_),
    .Y(_2321_));
 sky130_fd_sc_hd__a21oi_2 _6516_ (.A1(_2315_),
    .A2(_2320_),
    .B1(_2321_),
    .Y(_2322_));
 sky130_fd_sc_hd__a21o_1 _6517_ (.A1(_2295_),
    .A2(_2303_),
    .B1(_2322_),
    .X(_2323_));
 sky130_fd_sc_hd__a21o_1 _6518_ (.A1(_2173_),
    .A2(_2179_),
    .B1(_2181_),
    .X(_2324_));
 sky130_fd_sc_hd__nand3_1 _6519_ (.A(_2173_),
    .B(_2179_),
    .C(_2181_),
    .Y(_2325_));
 sky130_fd_sc_hd__nand2_1 _6520_ (.A(_2324_),
    .B(_2325_),
    .Y(_2326_));
 sky130_fd_sc_hd__nand2_1 _6521_ (.A(_2216_),
    .B(_2326_),
    .Y(_2328_));
 sky130_fd_sc_hd__nand2_1 _6522_ (.A(_2222_),
    .B(_2328_),
    .Y(_2329_));
 sky130_fd_sc_hd__nand3_1 _6523_ (.A(_2322_),
    .B(_2295_),
    .C(_2303_),
    .Y(_2330_));
 sky130_fd_sc_hd__nand3_1 _6524_ (.A(_2323_),
    .B(_2329_),
    .C(_2330_),
    .Y(_2331_));
 sky130_fd_sc_hd__a21boi_1 _6525_ (.A1(_2216_),
    .A2(_2326_),
    .B1_N(_2222_),
    .Y(_2332_));
 sky130_fd_sc_hd__nand2_1 _6526_ (.A(_2295_),
    .B(_2303_),
    .Y(_2333_));
 sky130_fd_sc_hd__nand2_1 _6527_ (.A(_2333_),
    .B(_2322_),
    .Y(_2334_));
 sky130_fd_sc_hd__inv_2 _6528_ (.A(_2320_),
    .Y(_2335_));
 sky130_fd_sc_hd__nand2_1 _6529_ (.A(_2312_),
    .B(_2314_),
    .Y(_2336_));
 sky130_fd_sc_hd__a21o_1 _6530_ (.A1(_2312_),
    .A2(_2320_),
    .B1(_2314_),
    .X(_2337_));
 sky130_fd_sc_hd__o21ai_2 _6531_ (.A1(_2335_),
    .A2(_2336_),
    .B1(_2337_),
    .Y(_2339_));
 sky130_fd_sc_hd__nand3_1 _6532_ (.A(_2339_),
    .B(_2295_),
    .C(_2303_),
    .Y(_2340_));
 sky130_fd_sc_hd__nand3_2 _6533_ (.A(_2332_),
    .B(_2334_),
    .C(_2340_),
    .Y(_2341_));
 sky130_fd_sc_hd__o211ai_1 _6534_ (.A1(_2264_),
    .A2(_2265_),
    .B1(_2331_),
    .C1(_2341_),
    .Y(_2342_));
 sky130_fd_sc_hd__nand2_1 _6535_ (.A(_2331_),
    .B(_2341_),
    .Y(_2343_));
 sky130_fd_sc_hd__nor2_1 _6536_ (.A(_2264_),
    .B(_2265_),
    .Y(_2344_));
 sky130_fd_sc_hd__nand2_1 _6537_ (.A(_2343_),
    .B(_2344_),
    .Y(_2345_));
 sky130_fd_sc_hd__nand3_1 _6538_ (.A(_2262_),
    .B(_2342_),
    .C(_2345_),
    .Y(_2346_));
 sky130_fd_sc_hd__o21ai_1 _6539_ (.A1(_2264_),
    .A2(_2265_),
    .B1(_2343_),
    .Y(_2347_));
 sky130_fd_sc_hd__and3_1 _6540_ (.A(_2322_),
    .B(_2295_),
    .C(_2303_),
    .X(_2348_));
 sky130_fd_sc_hd__nand2_1 _6541_ (.A(_2329_),
    .B(_2323_),
    .Y(_2350_));
 sky130_fd_sc_hd__o211ai_2 _6542_ (.A1(_2348_),
    .A2(_2350_),
    .B1(_2341_),
    .C1(_2344_),
    .Y(_2351_));
 sky130_fd_sc_hd__nand2_1 _6543_ (.A(_2233_),
    .B(_2237_),
    .Y(_2352_));
 sky130_fd_sc_hd__nand2_1 _6544_ (.A(_2228_),
    .B(_2352_),
    .Y(_2353_));
 sky130_fd_sc_hd__nand3_2 _6545_ (.A(_2347_),
    .B(_2351_),
    .C(_2353_),
    .Y(_2354_));
 sky130_fd_sc_hd__a21o_1 _6546_ (.A1(_2346_),
    .A2(_2354_),
    .B1(_2236_),
    .X(_2355_));
 sky130_fd_sc_hd__nand3_1 _6547_ (.A(_2346_),
    .B(_2354_),
    .C(_2236_),
    .Y(_2356_));
 sky130_fd_sc_hd__a32o_1 _6548_ (.A1(_2162_),
    .A2(_2238_),
    .A3(_2239_),
    .B1(_2245_),
    .B2(_2246_),
    .X(_2357_));
 sky130_fd_sc_hd__a21o_1 _6549_ (.A1(_2355_),
    .A2(_2356_),
    .B1(_2357_),
    .X(_2358_));
 sky130_fd_sc_hd__nand3_1 _6550_ (.A(_2357_),
    .B(_2355_),
    .C(_2356_),
    .Y(_2359_));
 sky130_fd_sc_hd__a21boi_1 _6551_ (.A1(_2260_),
    .A2(_2253_),
    .B1_N(_2255_),
    .Y(_2361_));
 sky130_fd_sc_hd__a21oi_1 _6552_ (.A1(_2358_),
    .A2(_2359_),
    .B1(_2361_),
    .Y(_2362_));
 sky130_fd_sc_hd__and3_1 _6553_ (.A(_2361_),
    .B(_2359_),
    .C(_2358_),
    .X(_2363_));
 sky130_fd_sc_hd__or2_1 _6554_ (.A(_2362_),
    .B(_2363_),
    .X(_2364_));
 sky130_fd_sc_hd__clkbuf_1 _6555_ (.A(_2364_),
    .X(_0092_));
 sky130_fd_sc_hd__nand2_1 _6556_ (.A(_2346_),
    .B(_2236_),
    .Y(_2365_));
 sky130_fd_sc_hd__a21boi_2 _6557_ (.A1(_2344_),
    .A2(_2341_),
    .B1_N(_2331_),
    .Y(_2366_));
 sky130_fd_sc_hd__and3_1 _6558_ (.A(_2336_),
    .B(_2234_),
    .C(_2320_),
    .X(_2367_));
 sky130_fd_sc_hd__o22a_2 _6559_ (.A1(_2013_),
    .A2(_2124_),
    .B1(_2335_),
    .B2(_2315_),
    .X(_2368_));
 sky130_fd_sc_hd__a21boi_1 _6560_ (.A1(_2322_),
    .A2(_2303_),
    .B1_N(_2295_),
    .Y(_2369_));
 sky130_fd_sc_hd__nand3_1 _6561_ (.A(net264),
    .B(net222),
    .C(net216),
    .Y(_2371_));
 sky130_fd_sc_hd__o21a_1 _6562_ (.A1(net222),
    .A2(net216),
    .B1(net264),
    .X(_2372_));
 sky130_fd_sc_hd__o2bb2ai_2 _6563_ (.A1_N(_2371_),
    .A2_N(_2372_),
    .B1(_1423_),
    .B2(_1366_),
    .Y(_2373_));
 sky130_fd_sc_hd__nand2_2 _6564_ (.A(net264),
    .B(net222),
    .Y(_2374_));
 sky130_fd_sc_hd__o211a_1 _6565_ (.A1(net223),
    .A2(net216),
    .B1(net263),
    .C1(net230),
    .X(_2375_));
 sky130_fd_sc_hd__o21ai_2 _6566_ (.A1(_1367_),
    .A2(_2374_),
    .B1(_2375_),
    .Y(_2376_));
 sky130_fd_sc_hd__a22oi_1 _6567_ (.A1(net303),
    .A2(net204),
    .B1(net314),
    .B2(net198),
    .Y(_2377_));
 sky130_fd_sc_hd__o21ai_1 _6568_ (.A1(_2299_),
    .A2(_2377_),
    .B1(_2284_),
    .Y(_2378_));
 sky130_fd_sc_hd__nand3_1 _6569_ (.A(_2373_),
    .B(_2376_),
    .C(_2378_),
    .Y(_2379_));
 sky130_fd_sc_hd__nand2_1 _6570_ (.A(net264),
    .B(net216),
    .Y(_2380_));
 sky130_fd_sc_hd__a21boi_4 _6571_ (.A1(_2374_),
    .A2(_2380_),
    .B1_N(_2371_),
    .Y(_2382_));
 sky130_fd_sc_hd__o211ai_4 _6572_ (.A1(_1367_),
    .A2(_2374_),
    .B1(_2372_),
    .C1(_1366_),
    .Y(_2383_));
 sky130_fd_sc_hd__o21a_1 _6573_ (.A1(_2299_),
    .A2(_2377_),
    .B1(_2282_),
    .X(_2384_));
 sky130_fd_sc_hd__o211ai_2 _6574_ (.A1(_2177_),
    .A2(_2382_),
    .B1(_2383_),
    .C1(_2384_),
    .Y(_2385_));
 sky130_fd_sc_hd__a21oi_2 _6575_ (.A1(_2177_),
    .A2(_2304_),
    .B1(_2307_),
    .Y(_2386_));
 sky130_fd_sc_hd__and3_1 _6576_ (.A(_2379_),
    .B(_2385_),
    .C(_2386_),
    .X(_2387_));
 sky130_fd_sc_hd__nand2_1 _6577_ (.A(_2379_),
    .B(_2385_),
    .Y(_2388_));
 sky130_fd_sc_hd__o311a_1 _6578_ (.A1(_3176_),
    .A2(_1332_),
    .A3(_2307_),
    .B1(_2304_),
    .C1(_2388_),
    .X(_2389_));
 sky130_fd_sc_hd__a22oi_2 _6579_ (.A1(net290),
    .A2(net204),
    .B1(net198),
    .B2(net303),
    .Y(_2390_));
 sky130_fd_sc_hd__nand2_1 _6580_ (.A(net279),
    .B(net212),
    .Y(_2391_));
 sky130_fd_sc_hd__a41o_1 _6581_ (.A1(net303),
    .A2(net290),
    .A3(net204),
    .A4(net198),
    .B1(_2391_),
    .X(_2393_));
 sky130_fd_sc_hd__a22o_1 _6582_ (.A1(net290),
    .A2(net205),
    .B1(net199),
    .B2(net303),
    .X(_2394_));
 sky130_fd_sc_hd__nand4_1 _6583_ (.A(net303),
    .B(net290),
    .C(net205),
    .D(net199),
    .Y(_2395_));
 sky130_fd_sc_hd__a22o_1 _6584_ (.A1(net279),
    .A2(net212),
    .B1(_2394_),
    .B2(_2395_),
    .X(_2396_));
 sky130_fd_sc_hd__o21ai_2 _6585_ (.A1(_2390_),
    .A2(_2393_),
    .B1(_2396_),
    .Y(_2397_));
 sky130_fd_sc_hd__o2bb2ai_4 _6586_ (.A1_N(net326),
    .A2_N(net186),
    .B1(net338),
    .B2(_1953_),
    .Y(_2398_));
 sky130_fd_sc_hd__nand4b_4 _6587_ (.A_N(net338),
    .B(net326),
    .C(net184),
    .D(net179),
    .Y(_2399_));
 sky130_fd_sc_hd__nand2_1 _6588_ (.A(net313),
    .B(net192),
    .Y(_2400_));
 sky130_fd_sc_hd__a21oi_4 _6589_ (.A1(_2398_),
    .A2(_2399_),
    .B1(_2400_),
    .Y(_2401_));
 sky130_fd_sc_hd__a22oi_4 _6590_ (.A1(net326),
    .A2(net186),
    .B1(_2120_),
    .B2(net180),
    .Y(_2402_));
 sky130_fd_sc_hd__o21ai_4 _6591_ (.A1(_2848_),
    .A2(_1642_),
    .B1(_2399_),
    .Y(_2404_));
 sky130_fd_sc_hd__o221ai_4 _6592_ (.A1(_2277_),
    .A2(_2271_),
    .B1(_2402_),
    .B2(_2404_),
    .C1(_2269_),
    .Y(_2405_));
 sky130_fd_sc_hd__and4b_1 _6593_ (.A_N(net338),
    .B(net326),
    .C(net186),
    .D(net180),
    .X(_2406_));
 sky130_fd_sc_hd__o22ai_1 _6594_ (.A1(_2973_),
    .A2(_2199_),
    .B1(_2402_),
    .B2(_2406_),
    .Y(_2407_));
 sky130_fd_sc_hd__o21ai_1 _6595_ (.A1(_2277_),
    .A2(_2271_),
    .B1(_2269_),
    .Y(_2408_));
 sky130_fd_sc_hd__nand4_1 _6596_ (.A(_2398_),
    .B(_2399_),
    .C(net313),
    .D(net192),
    .Y(_2409_));
 sky130_fd_sc_hd__nand3_2 _6597_ (.A(_2407_),
    .B(_2408_),
    .C(_2409_),
    .Y(_2410_));
 sky130_fd_sc_hd__o21ai_1 _6598_ (.A1(_2401_),
    .A2(_2405_),
    .B1(_2410_),
    .Y(_2411_));
 sky130_fd_sc_hd__nand2_1 _6599_ (.A(_2397_),
    .B(_2411_),
    .Y(_2412_));
 sky130_fd_sc_hd__nand2_1 _6600_ (.A(_2268_),
    .B(_2269_),
    .Y(_2413_));
 sky130_fd_sc_hd__a22oi_2 _6601_ (.A1(_2192_),
    .A2(_2266_),
    .B1(_2413_),
    .B2(_2274_),
    .Y(_2415_));
 sky130_fd_sc_hd__nand2_1 _6602_ (.A(_2291_),
    .B(_2292_),
    .Y(_2416_));
 sky130_fd_sc_hd__a22oi_2 _6603_ (.A1(_2270_),
    .A2(_2415_),
    .B1(_2281_),
    .B2(_2416_),
    .Y(_2417_));
 sky130_fd_sc_hd__o21a_1 _6604_ (.A1(_2390_),
    .A2(_2393_),
    .B1(_2396_),
    .X(_2418_));
 sky130_fd_sc_hd__o211ai_2 _6605_ (.A1(_2401_),
    .A2(_2405_),
    .B1(_2410_),
    .C1(_2418_),
    .Y(_2419_));
 sky130_fd_sc_hd__nand3_2 _6606_ (.A(_2412_),
    .B(_2417_),
    .C(_2419_),
    .Y(_2420_));
 sky130_fd_sc_hd__a22o_1 _6607_ (.A1(_2270_),
    .A2(_2415_),
    .B1(_2281_),
    .B2(_2416_),
    .X(_2421_));
 sky130_fd_sc_hd__o211ai_1 _6608_ (.A1(_2401_),
    .A2(_2405_),
    .B1(_2397_),
    .C1(_2410_),
    .Y(_2422_));
 sky130_fd_sc_hd__nand2_1 _6609_ (.A(_2411_),
    .B(_2418_),
    .Y(_2423_));
 sky130_fd_sc_hd__nand3_2 _6610_ (.A(_2421_),
    .B(_2422_),
    .C(_2423_),
    .Y(_2424_));
 sky130_fd_sc_hd__o211ai_1 _6611_ (.A1(_2387_),
    .A2(_2389_),
    .B1(_2420_),
    .C1(_2424_),
    .Y(_2426_));
 sky130_fd_sc_hd__nand2_1 _6612_ (.A(_2388_),
    .B(_2386_),
    .Y(_2427_));
 sky130_fd_sc_hd__inv_2 _6613_ (.A(_2427_),
    .Y(_2428_));
 sky130_fd_sc_hd__a21oi_1 _6614_ (.A1(_2310_),
    .A2(_2306_),
    .B1(_2388_),
    .Y(_2429_));
 sky130_fd_sc_hd__o2bb2ai_1 _6615_ (.A1_N(_2420_),
    .A2_N(_2424_),
    .B1(_2428_),
    .B2(_2429_),
    .Y(_2430_));
 sky130_fd_sc_hd__nand3_2 _6616_ (.A(_2369_),
    .B(_2426_),
    .C(_2430_),
    .Y(_2431_));
 sky130_fd_sc_hd__nand2_1 _6617_ (.A(_2276_),
    .B(_2281_),
    .Y(_2432_));
 sky130_fd_sc_hd__a21oi_1 _6618_ (.A1(_2432_),
    .A2(_2288_),
    .B1(_2290_),
    .Y(_2433_));
 sky130_fd_sc_hd__a31o_1 _6619_ (.A1(_2267_),
    .A2(_2270_),
    .A3(_2275_),
    .B1(_2296_),
    .X(_2434_));
 sky130_fd_sc_hd__a22oi_2 _6620_ (.A1(_2433_),
    .A2(_2434_),
    .B1(_2339_),
    .B2(_2295_),
    .Y(_2435_));
 sky130_fd_sc_hd__o211ai_1 _6621_ (.A1(_2428_),
    .A2(_2429_),
    .B1(_2420_),
    .C1(_2424_),
    .Y(_2437_));
 sky130_fd_sc_hd__o2bb2ai_1 _6622_ (.A1_N(_2420_),
    .A2_N(_2424_),
    .B1(_2387_),
    .B2(_2389_),
    .Y(_2438_));
 sky130_fd_sc_hd__nand3_2 _6623_ (.A(_2435_),
    .B(_2437_),
    .C(_2438_),
    .Y(_2439_));
 sky130_fd_sc_hd__o211ai_2 _6624_ (.A1(_2367_),
    .A2(_2368_),
    .B1(_2431_),
    .C1(_2439_),
    .Y(_2440_));
 sky130_fd_sc_hd__nand2_1 _6625_ (.A(_2431_),
    .B(_2439_),
    .Y(_2441_));
 sky130_fd_sc_hd__nor2_1 _6626_ (.A(_2367_),
    .B(_2368_),
    .Y(_2442_));
 sky130_fd_sc_hd__nand2_1 _6627_ (.A(_2441_),
    .B(_2442_),
    .Y(_2443_));
 sky130_fd_sc_hd__nand3_1 _6628_ (.A(_2366_),
    .B(_2440_),
    .C(_2443_),
    .Y(_2444_));
 sky130_fd_sc_hd__o2bb2ai_1 _6629_ (.A1_N(_2344_),
    .A2_N(_2341_),
    .B1(_2348_),
    .B2(_2350_),
    .Y(_2445_));
 sky130_fd_sc_hd__o2bb2ai_1 _6630_ (.A1_N(_2431_),
    .A2_N(_2439_),
    .B1(_2367_),
    .B2(_2368_),
    .Y(_2446_));
 sky130_fd_sc_hd__nand3_1 _6631_ (.A(_2431_),
    .B(_2439_),
    .C(_2442_),
    .Y(_2448_));
 sky130_fd_sc_hd__nand3_2 _6632_ (.A(_2445_),
    .B(_2446_),
    .C(_2448_),
    .Y(_2449_));
 sky130_fd_sc_hd__o21ai_2 _6633_ (.A1(_2013_),
    .A2(_2124_),
    .B1(_2263_),
    .Y(_2450_));
 sky130_fd_sc_hd__a21o_1 _6634_ (.A1(_2444_),
    .A2(_2449_),
    .B1(_2450_),
    .X(_2451_));
 sky130_fd_sc_hd__nand3_2 _6635_ (.A(_2450_),
    .B(_2444_),
    .C(_2449_),
    .Y(_2452_));
 sky130_fd_sc_hd__a22oi_4 _6636_ (.A1(_2354_),
    .A2(_2365_),
    .B1(_2451_),
    .B2(_2452_),
    .Y(_2453_));
 sky130_fd_sc_hd__and3_1 _6637_ (.A(_2262_),
    .B(_2342_),
    .C(_2345_),
    .X(_2454_));
 sky130_fd_sc_hd__a31oi_1 _6638_ (.A1(_2347_),
    .A2(_2351_),
    .A3(_2353_),
    .B1(_2236_),
    .Y(_2455_));
 sky130_fd_sc_hd__o211a_1 _6639_ (.A1(_2454_),
    .A2(_2455_),
    .B1(_2451_),
    .C1(_2452_),
    .X(_2456_));
 sky130_fd_sc_hd__nor2_1 _6640_ (.A(_2453_),
    .B(_2456_),
    .Y(_2457_));
 sky130_fd_sc_hd__nand2_1 _6641_ (.A(_2255_),
    .B(_2359_),
    .Y(_2459_));
 sky130_fd_sc_hd__a22oi_2 _6642_ (.A1(_2156_),
    .A2(_2257_),
    .B1(_2358_),
    .B2(_2459_),
    .Y(_2460_));
 sky130_fd_sc_hd__o21ai_2 _6643_ (.A1(_2050_),
    .A2(_2259_),
    .B1(_2460_),
    .Y(_2461_));
 sky130_fd_sc_hd__a21bo_1 _6644_ (.A1(_2253_),
    .A2(_2358_),
    .B1_N(_2359_),
    .X(_2462_));
 sky130_fd_sc_hd__nand2_1 _6645_ (.A(_2461_),
    .B(_2462_),
    .Y(_2463_));
 sky130_fd_sc_hd__xnor2_1 _6646_ (.A(_2457_),
    .B(_2463_),
    .Y(_0093_));
 sky130_fd_sc_hd__a2bb2o_1 _6647_ (.A1_N(_2013_),
    .A2_N(_2124_),
    .B1(_2320_),
    .B2(_2336_),
    .X(_2464_));
 sky130_fd_sc_hd__a21oi_1 _6648_ (.A1(_2395_),
    .A2(_2391_),
    .B1(_2390_),
    .Y(_2465_));
 sky130_fd_sc_hd__a21o_1 _6649_ (.A1(_2373_),
    .A2(_2376_),
    .B1(_2465_),
    .X(_2466_));
 sky130_fd_sc_hd__a31o_1 _6650_ (.A1(net263),
    .A2(net222),
    .A3(net216),
    .B1(_2375_),
    .X(_2467_));
 sky130_fd_sc_hd__buf_4 _6651_ (.A(_2373_),
    .X(_2469_));
 sky130_fd_sc_hd__buf_6 _6652_ (.A(_2376_),
    .X(_2470_));
 sky130_fd_sc_hd__nand3_2 _6653_ (.A(_2469_),
    .B(_2470_),
    .C(_2465_),
    .Y(_2471_));
 sky130_fd_sc_hd__and3_1 _6654_ (.A(_2466_),
    .B(_2467_),
    .C(_2471_),
    .X(_2472_));
 sky130_fd_sc_hd__buf_2 _6655_ (.A(_2467_),
    .X(_2473_));
 sky130_fd_sc_hd__a21oi_2 _6656_ (.A1(_2471_),
    .A2(_2466_),
    .B1(_2473_),
    .Y(_2474_));
 sky130_fd_sc_hd__o2bb2ai_4 _6657_ (.A1_N(net313),
    .A2_N(net185),
    .B1(net326),
    .B2(_1953_),
    .Y(_2475_));
 sky130_fd_sc_hd__nand4_2 _6658_ (.A(_1782_),
    .B(net313),
    .C(net185),
    .D(net180),
    .Y(_2476_));
 sky130_fd_sc_hd__a22oi_2 _6659_ (.A1(net302),
    .A2(net192),
    .B1(_2475_),
    .B2(_2476_),
    .Y(_2477_));
 sky130_fd_sc_hd__nand3b_2 _6660_ (.A_N(net321),
    .B(net313),
    .C(net185),
    .Y(_2478_));
 sky130_fd_sc_hd__o2111a_1 _6661_ (.A1(_1958_),
    .A2(_2478_),
    .B1(net302),
    .C1(net194),
    .D1(_2475_),
    .X(_2480_));
 sky130_fd_sc_hd__o2bb2ai_4 _6662_ (.A1_N(_2398_),
    .A2_N(_2404_),
    .B1(_2477_),
    .B2(_2480_),
    .Y(_2481_));
 sky130_fd_sc_hd__nor2_1 _6663_ (.A(_2400_),
    .B(_2402_),
    .Y(_2482_));
 sky130_fd_sc_hd__o2111ai_4 _6664_ (.A1(_1958_),
    .A2(_2478_),
    .B1(net302),
    .C1(net194),
    .D1(_2475_),
    .Y(_2483_));
 sky130_fd_sc_hd__o2bb2ai_2 _6665_ (.A1_N(_2475_),
    .A2_N(_2476_),
    .B1(_3022_),
    .B2(_2199_),
    .Y(_2484_));
 sky130_fd_sc_hd__o211ai_4 _6666_ (.A1(_2406_),
    .A2(_2482_),
    .B1(_2483_),
    .C1(_2484_),
    .Y(_2485_));
 sky130_fd_sc_hd__a22oi_2 _6667_ (.A1(net279),
    .A2(net203),
    .B1(net197),
    .B2(net290),
    .Y(_2486_));
 sky130_fd_sc_hd__nand2_2 _6668_ (.A(net267),
    .B(net212),
    .Y(_2487_));
 sky130_fd_sc_hd__a41o_1 _6669_ (.A1(net291),
    .A2(net279),
    .A3(net203),
    .A4(net197),
    .B1(_2487_),
    .X(_2488_));
 sky130_fd_sc_hd__nand4_1 _6670_ (.A(net291),
    .B(net279),
    .C(net203),
    .D(net197),
    .Y(_2489_));
 sky130_fd_sc_hd__nand2_1 _6671_ (.A(net291),
    .B(net197),
    .Y(_2491_));
 sky130_fd_sc_hd__nand2_1 _6672_ (.A(net279),
    .B(net203),
    .Y(_2492_));
 sky130_fd_sc_hd__nand2_1 _6673_ (.A(_2491_),
    .B(_2492_),
    .Y(_2493_));
 sky130_fd_sc_hd__a22o_1 _6674_ (.A1(net266),
    .A2(net212),
    .B1(_2489_),
    .B2(_2493_),
    .X(_2494_));
 sky130_fd_sc_hd__o21a_1 _6675_ (.A1(_2486_),
    .A2(_2488_),
    .B1(_2494_),
    .X(_2495_));
 sky130_fd_sc_hd__a21oi_2 _6676_ (.A1(_2481_),
    .A2(_2485_),
    .B1(_2495_),
    .Y(_2496_));
 sky130_fd_sc_hd__nand2_1 _6677_ (.A(_2410_),
    .B(_2397_),
    .Y(_2497_));
 sky130_fd_sc_hd__nand3_1 _6678_ (.A(_2481_),
    .B(_2485_),
    .C(_2495_),
    .Y(_2498_));
 sky130_fd_sc_hd__o211ai_4 _6679_ (.A1(_2401_),
    .A2(_2405_),
    .B1(_2497_),
    .C1(_2498_),
    .Y(_2499_));
 sky130_fd_sc_hd__a22oi_2 _6680_ (.A1(_2398_),
    .A2(_2404_),
    .B1(_2484_),
    .B2(_2483_),
    .Y(_2500_));
 sky130_fd_sc_hd__o211a_1 _6681_ (.A1(_2406_),
    .A2(_2482_),
    .B1(_2483_),
    .C1(_2484_),
    .X(_2502_));
 sky130_fd_sc_hd__o21ai_1 _6682_ (.A1(_2500_),
    .A2(_2502_),
    .B1(_2495_),
    .Y(_2503_));
 sky130_fd_sc_hd__o21ai_1 _6683_ (.A1(_2401_),
    .A2(_2405_),
    .B1(_2497_),
    .Y(_2504_));
 sky130_fd_sc_hd__o21ai_2 _6684_ (.A1(_2486_),
    .A2(_2488_),
    .B1(_2494_),
    .Y(_2505_));
 sky130_fd_sc_hd__nand3_1 _6685_ (.A(_2481_),
    .B(_2485_),
    .C(_2505_),
    .Y(_2506_));
 sky130_fd_sc_hd__nand3_4 _6686_ (.A(_2503_),
    .B(_2504_),
    .C(_2506_),
    .Y(_2507_));
 sky130_fd_sc_hd__o221ai_4 _6687_ (.A1(_2472_),
    .A2(_2474_),
    .B1(_2496_),
    .B2(_2499_),
    .C1(_2507_),
    .Y(_2508_));
 sky130_fd_sc_hd__o21ai_1 _6688_ (.A1(_2496_),
    .A2(_2499_),
    .B1(_2507_),
    .Y(_2509_));
 sky130_fd_sc_hd__nor2_1 _6689_ (.A(_2472_),
    .B(_2474_),
    .Y(_2510_));
 sky130_fd_sc_hd__nand2_1 _6690_ (.A(_2509_),
    .B(_2510_),
    .Y(_2511_));
 sky130_fd_sc_hd__nand3b_1 _6691_ (.A_N(_2386_),
    .B(_2385_),
    .C(_2379_),
    .Y(_2513_));
 sky130_fd_sc_hd__nand2_1 _6692_ (.A(_2427_),
    .B(_2513_),
    .Y(_2514_));
 sky130_fd_sc_hd__a21oi_1 _6693_ (.A1(_2397_),
    .A2(_2411_),
    .B1(_2421_),
    .Y(_2515_));
 sky130_fd_sc_hd__a22oi_2 _6694_ (.A1(_2514_),
    .A2(_2424_),
    .B1(_2515_),
    .B2(_2419_),
    .Y(_2516_));
 sky130_fd_sc_hd__nand3_2 _6695_ (.A(_2508_),
    .B(_2511_),
    .C(_2516_),
    .Y(_2517_));
 sky130_fd_sc_hd__o21ai_1 _6696_ (.A1(_2472_),
    .A2(_2474_),
    .B1(_2509_),
    .Y(_2518_));
 sky130_fd_sc_hd__o211ai_1 _6697_ (.A1(_2496_),
    .A2(_2499_),
    .B1(_2507_),
    .C1(_2510_),
    .Y(_2519_));
 sky130_fd_sc_hd__nand2_1 _6698_ (.A(_2424_),
    .B(_2514_),
    .Y(_2520_));
 sky130_fd_sc_hd__nand2_1 _6699_ (.A(_2420_),
    .B(_2520_),
    .Y(_2521_));
 sky130_fd_sc_hd__nand3_2 _6700_ (.A(_2518_),
    .B(_2519_),
    .C(_2521_),
    .Y(_2522_));
 sky130_fd_sc_hd__clkbuf_4 _6701_ (.A(_2234_),
    .X(_2524_));
 sky130_fd_sc_hd__a32oi_2 _6702_ (.A1(_2378_),
    .A2(_2469_),
    .A3(_2470_),
    .B1(_2385_),
    .B2(_2386_),
    .Y(_2525_));
 sky130_fd_sc_hd__nor2_1 _6703_ (.A(_2524_),
    .B(_2525_),
    .Y(_2526_));
 sky130_fd_sc_hd__and2_1 _6704_ (.A(_2234_),
    .B(_2525_),
    .X(_2527_));
 sky130_fd_sc_hd__or2_1 _6705_ (.A(_2526_),
    .B(_2527_),
    .X(_2528_));
 sky130_fd_sc_hd__a21oi_2 _6706_ (.A1(_2517_),
    .A2(_2522_),
    .B1(_2528_),
    .Y(_2529_));
 sky130_fd_sc_hd__nand2_1 _6707_ (.A(_2431_),
    .B(_2442_),
    .Y(_2530_));
 sky130_fd_sc_hd__nand3_1 _6708_ (.A(_2517_),
    .B(_2522_),
    .C(_2528_),
    .Y(_2531_));
 sky130_fd_sc_hd__nand3_2 _6709_ (.A(_2439_),
    .B(_2530_),
    .C(_2531_),
    .Y(_2532_));
 sky130_fd_sc_hd__o2bb2ai_1 _6710_ (.A1_N(_2517_),
    .A2_N(_2522_),
    .B1(_2526_),
    .B2(_2527_),
    .Y(_2533_));
 sky130_fd_sc_hd__nand2_1 _6711_ (.A(_2439_),
    .B(_2530_),
    .Y(_2535_));
 sky130_fd_sc_hd__nand3b_1 _6712_ (.A_N(_2528_),
    .B(_2522_),
    .C(_2517_),
    .Y(_2536_));
 sky130_fd_sc_hd__nand3_1 _6713_ (.A(_2533_),
    .B(_2535_),
    .C(_2536_),
    .Y(_2537_));
 sky130_fd_sc_hd__o21ai_1 _6714_ (.A1(_2529_),
    .A2(_2532_),
    .B1(_2537_),
    .Y(_2538_));
 sky130_fd_sc_hd__nand2_1 _6715_ (.A(_2464_),
    .B(_2538_),
    .Y(_2539_));
 sky130_fd_sc_hd__o211ai_2 _6716_ (.A1(_2529_),
    .A2(_2532_),
    .B1(_2537_),
    .C1(_2368_),
    .Y(_2540_));
 sky130_fd_sc_hd__a32oi_4 _6717_ (.A1(_2366_),
    .A2(_2440_),
    .A3(_2443_),
    .B1(_2449_),
    .B2(_2450_),
    .Y(_2541_));
 sky130_fd_sc_hd__nand3_1 _6718_ (.A(_2539_),
    .B(_2540_),
    .C(_2541_),
    .Y(_2542_));
 sky130_fd_sc_hd__nand2_1 _6719_ (.A(_2538_),
    .B(_2368_),
    .Y(_2543_));
 sky130_fd_sc_hd__o211ai_1 _6720_ (.A1(_2529_),
    .A2(_2532_),
    .B1(_2537_),
    .C1(_2464_),
    .Y(_2544_));
 sky130_fd_sc_hd__a21boi_1 _6721_ (.A1(_2444_),
    .A2(_2264_),
    .B1_N(_2449_),
    .Y(_2546_));
 sky130_fd_sc_hd__nand3_1 _6722_ (.A(_2543_),
    .B(_2544_),
    .C(_2546_),
    .Y(_2547_));
 sky130_fd_sc_hd__and2_1 _6723_ (.A(_2542_),
    .B(_2547_),
    .X(_2548_));
 sky130_fd_sc_hd__a31oi_1 _6724_ (.A1(_2461_),
    .A2(_2462_),
    .A3(_2457_),
    .B1(_2453_),
    .Y(_2549_));
 sky130_fd_sc_hd__xnor2_1 _6725_ (.A(_2548_),
    .B(_2549_),
    .Y(_0094_));
 sky130_fd_sc_hd__nand3_1 _6726_ (.A(_2250_),
    .B(_2252_),
    .C(_2359_),
    .Y(_2550_));
 sky130_fd_sc_hd__and4_1 _6727_ (.A(_2457_),
    .B(_2548_),
    .C(_2550_),
    .D(_2358_),
    .X(_2551_));
 sky130_fd_sc_hd__a32oi_4 _6728_ (.A1(_2539_),
    .A2(_2540_),
    .A3(_2541_),
    .B1(_2453_),
    .B2(_2547_),
    .Y(_2552_));
 sky130_fd_sc_hd__a21boi_1 _6729_ (.A1(_2461_),
    .A2(_2551_),
    .B1_N(_2552_),
    .Y(_2553_));
 sky130_fd_sc_hd__nand2_1 _6730_ (.A(_2508_),
    .B(_2511_),
    .Y(_2554_));
 sky130_fd_sc_hd__nand2_1 _6731_ (.A(_2522_),
    .B(_2528_),
    .Y(_2556_));
 sky130_fd_sc_hd__o21ai_1 _6732_ (.A1(_2554_),
    .A2(_2521_),
    .B1(_2556_),
    .Y(_2557_));
 sky130_fd_sc_hd__nand4_4 _6733_ (.A(_2794_),
    .B(net185),
    .C(net180),
    .D(net304),
    .Y(_2558_));
 sky130_fd_sc_hd__o2bb2ai_2 _6734_ (.A1_N(net302),
    .A2_N(net185),
    .B1(net315),
    .B2(_1953_),
    .Y(_2559_));
 sky130_fd_sc_hd__o2bb2ai_2 _6735_ (.A1_N(_2558_),
    .A2_N(_2559_),
    .B1(_0509_),
    .B2(_1643_),
    .Y(_2560_));
 sky130_fd_sc_hd__nor2_1 _6736_ (.A(_3381_),
    .B(_1641_),
    .Y(_2561_));
 sky130_fd_sc_hd__nand3_2 _6737_ (.A(_2559_),
    .B(_2561_),
    .C(_2558_),
    .Y(_2562_));
 sky130_fd_sc_hd__nand2_1 _6738_ (.A(net302),
    .B(net192),
    .Y(_2563_));
 sky130_fd_sc_hd__a22oi_2 _6739_ (.A1(net313),
    .A2(net185),
    .B1(_2886_),
    .B2(net180),
    .Y(_2564_));
 sky130_fd_sc_hd__o21ai_2 _6740_ (.A1(_2563_),
    .A2(_2564_),
    .B1(_2476_),
    .Y(_2565_));
 sky130_fd_sc_hd__a21oi_2 _6741_ (.A1(_2560_),
    .A2(_2562_),
    .B1(_2565_),
    .Y(_2567_));
 sky130_fd_sc_hd__and3_2 _6742_ (.A(_2565_),
    .B(_2560_),
    .C(_2562_),
    .X(_2568_));
 sky130_fd_sc_hd__nand4_2 _6743_ (.A(net279),
    .B(net267),
    .C(net205),
    .D(net199),
    .Y(_2569_));
 sky130_fd_sc_hd__nand2_1 _6744_ (.A(net279),
    .B(net199),
    .Y(_2570_));
 sky130_fd_sc_hd__nand2_1 _6745_ (.A(net267),
    .B(net205),
    .Y(_2571_));
 sky130_fd_sc_hd__nand2_1 _6746_ (.A(_2570_),
    .B(_2571_),
    .Y(_2572_));
 sky130_fd_sc_hd__and3_1 _6747_ (.A(_2487_),
    .B(_2569_),
    .C(_2572_),
    .X(_2573_));
 sky130_fd_sc_hd__a21oi_1 _6748_ (.A1(_2569_),
    .A2(_2572_),
    .B1(_2487_),
    .Y(_2574_));
 sky130_fd_sc_hd__nor2_1 _6749_ (.A(_2573_),
    .B(_2574_),
    .Y(_2575_));
 sky130_fd_sc_hd__o21ai_1 _6750_ (.A1(_2567_),
    .A2(_2568_),
    .B1(_2575_),
    .Y(_2576_));
 sky130_fd_sc_hd__o21ai_1 _6751_ (.A1(_2500_),
    .A2(_2505_),
    .B1(_2485_),
    .Y(_2578_));
 sky130_fd_sc_hd__a21o_1 _6752_ (.A1(_2560_),
    .A2(_2562_),
    .B1(_2565_),
    .X(_2579_));
 sky130_fd_sc_hd__nand3_2 _6753_ (.A(_2565_),
    .B(_2560_),
    .C(_2562_),
    .Y(_2580_));
 sky130_fd_sc_hd__o211ai_2 _6754_ (.A1(_2573_),
    .A2(_2574_),
    .B1(_2579_),
    .C1(_2580_),
    .Y(_2581_));
 sky130_fd_sc_hd__nand3_4 _6755_ (.A(_2576_),
    .B(_2578_),
    .C(_2581_),
    .Y(_2582_));
 sky130_fd_sc_hd__o2bb2a_1 _6756_ (.A1_N(_2569_),
    .A2_N(_2572_),
    .B1(_3058_),
    .B2(_1394_),
    .X(_2583_));
 sky130_fd_sc_hd__nor2_1 _6757_ (.A(_3342_),
    .B(_1394_),
    .Y(_2584_));
 sky130_fd_sc_hd__and3_1 _6758_ (.A(_2584_),
    .B(_2569_),
    .C(_2572_),
    .X(_2585_));
 sky130_fd_sc_hd__o211ai_2 _6759_ (.A1(_2583_),
    .A2(_2585_),
    .B1(_2579_),
    .C1(_2580_),
    .Y(_2586_));
 sky130_fd_sc_hd__nor2_1 _6760_ (.A(_2583_),
    .B(_2585_),
    .Y(_2587_));
 sky130_fd_sc_hd__o21ai_1 _6761_ (.A1(_2567_),
    .A2(_2568_),
    .B1(_2587_),
    .Y(_2589_));
 sky130_fd_sc_hd__a21oi_1 _6762_ (.A1(_2481_),
    .A2(_2495_),
    .B1(_2502_),
    .Y(_2590_));
 sky130_fd_sc_hd__nand3_2 _6763_ (.A(_2586_),
    .B(_2589_),
    .C(_2590_),
    .Y(_2591_));
 sky130_fd_sc_hd__o21ai_1 _6764_ (.A1(_2491_),
    .A2(_2492_),
    .B1(_2487_),
    .Y(_2592_));
 sky130_fd_sc_hd__nand4_2 _6765_ (.A(_2469_),
    .B(_2470_),
    .C(_2493_),
    .D(_2592_),
    .Y(_2593_));
 sky130_fd_sc_hd__o21a_1 _6766_ (.A1(_2487_),
    .A2(_2486_),
    .B1(_2489_),
    .X(_2594_));
 sky130_fd_sc_hd__o211ai_2 _6767_ (.A1(_2177_),
    .A2(_2382_),
    .B1(_2383_),
    .C1(_2594_),
    .Y(_2595_));
 sky130_fd_sc_hd__a21oi_1 _6768_ (.A1(_2593_),
    .A2(_2595_),
    .B1(_2467_),
    .Y(_2596_));
 sky130_fd_sc_hd__and3_1 _6769_ (.A(_2595_),
    .B(_2467_),
    .C(_2593_),
    .X(_2597_));
 sky130_fd_sc_hd__nor2_1 _6770_ (.A(_2596_),
    .B(_2597_),
    .Y(_2598_));
 sky130_fd_sc_hd__a21oi_2 _6771_ (.A1(_2582_),
    .A2(_2591_),
    .B1(_2598_),
    .Y(_2600_));
 sky130_fd_sc_hd__nor2_1 _6772_ (.A(_2496_),
    .B(_2499_),
    .Y(_2601_));
 sky130_fd_sc_hd__nand3_1 _6773_ (.A(_2582_),
    .B(_2591_),
    .C(_2598_),
    .Y(_2602_));
 sky130_fd_sc_hd__o211ai_2 _6774_ (.A1(_2510_),
    .A2(_2601_),
    .B1(_2602_),
    .C1(_2507_),
    .Y(_2603_));
 sky130_fd_sc_hd__nand3_1 _6775_ (.A(_2595_),
    .B(_2467_),
    .C(_2593_),
    .Y(_2604_));
 sky130_fd_sc_hd__nand2b_1 _6776_ (.A_N(_2596_),
    .B(_2604_),
    .Y(_2605_));
 sky130_fd_sc_hd__a21o_1 _6777_ (.A1(_2582_),
    .A2(_2591_),
    .B1(_2605_),
    .X(_2606_));
 sky130_fd_sc_hd__o21ai_1 _6778_ (.A1(_2510_),
    .A2(_2601_),
    .B1(_2507_),
    .Y(_2607_));
 sky130_fd_sc_hd__o211ai_1 _6779_ (.A1(_2596_),
    .A2(_2597_),
    .B1(_2582_),
    .C1(_2591_),
    .Y(_2608_));
 sky130_fd_sc_hd__nand3_1 _6780_ (.A(_2606_),
    .B(_2607_),
    .C(_2608_),
    .Y(_2609_));
 sky130_fd_sc_hd__nand3_1 _6781_ (.A(_2466_),
    .B(_2473_),
    .C(_2471_),
    .Y(_2611_));
 sky130_fd_sc_hd__and3_1 _6782_ (.A(_2611_),
    .B(_2524_),
    .C(_2471_),
    .X(_2612_));
 sky130_fd_sc_hd__a21oi_2 _6783_ (.A1(_2471_),
    .A2(_2611_),
    .B1(_2524_),
    .Y(_2613_));
 sky130_fd_sc_hd__nor2_1 _6784_ (.A(_2612_),
    .B(_2613_),
    .Y(_2614_));
 sky130_fd_sc_hd__o211ai_1 _6785_ (.A1(_2600_),
    .A2(_2603_),
    .B1(_2609_),
    .C1(_2614_),
    .Y(_2615_));
 sky130_fd_sc_hd__o21ai_1 _6786_ (.A1(_2600_),
    .A2(_2603_),
    .B1(_2609_),
    .Y(_2616_));
 sky130_fd_sc_hd__o21ai_1 _6787_ (.A1(_2612_),
    .A2(_2613_),
    .B1(_2616_),
    .Y(_2617_));
 sky130_fd_sc_hd__nand3b_1 _6788_ (.A_N(_2557_),
    .B(_2615_),
    .C(_2617_),
    .Y(_2618_));
 sky130_fd_sc_hd__nand2_1 _6789_ (.A(_2616_),
    .B(_2614_),
    .Y(_2619_));
 sky130_fd_sc_hd__o221ai_1 _6790_ (.A1(_2612_),
    .A2(_2613_),
    .B1(_2600_),
    .B2(_2603_),
    .C1(_2609_),
    .Y(_2620_));
 sky130_fd_sc_hd__nand3_1 _6791_ (.A(_2557_),
    .B(_2619_),
    .C(_2620_),
    .Y(_2622_));
 sky130_fd_sc_hd__a21o_1 _6792_ (.A1(_2618_),
    .A2(_2622_),
    .B1(_2526_),
    .X(_2623_));
 sky130_fd_sc_hd__nand3_1 _6793_ (.A(_2618_),
    .B(_2622_),
    .C(_2526_),
    .Y(_2624_));
 sky130_fd_sc_hd__o2bb2a_1 _6794_ (.A1_N(_2464_),
    .A2_N(_2537_),
    .B1(_2532_),
    .B2(_2529_),
    .X(_2625_));
 sky130_fd_sc_hd__a21o_1 _6795_ (.A1(_2623_),
    .A2(_2624_),
    .B1(_2625_),
    .X(_2626_));
 sky130_fd_sc_hd__nand3_1 _6796_ (.A(_2623_),
    .B(_2624_),
    .C(_2625_),
    .Y(_2627_));
 sky130_fd_sc_hd__nand2_2 _6797_ (.A(_2626_),
    .B(_2627_),
    .Y(_2628_));
 sky130_fd_sc_hd__xor2_1 _6798_ (.A(_2553_),
    .B(_2628_),
    .X(_0095_));
 sky130_fd_sc_hd__o21ai_1 _6799_ (.A1(_2628_),
    .A2(_2553_),
    .B1(_2627_),
    .Y(_2629_));
 sky130_fd_sc_hd__a2bb2oi_1 _6800_ (.A1_N(_2600_),
    .A2_N(_2603_),
    .B1(_2614_),
    .B2(_2609_),
    .Y(_2630_));
 sky130_fd_sc_hd__and3_1 _6801_ (.A(_2604_),
    .B(_2524_),
    .C(_2593_),
    .X(_2632_));
 sky130_fd_sc_hd__a21oi_2 _6802_ (.A1(_2593_),
    .A2(_2604_),
    .B1(_2524_),
    .Y(_2633_));
 sky130_fd_sc_hd__a21boi_2 _6803_ (.A1(_2487_),
    .A2(_2569_),
    .B1_N(_2572_),
    .Y(_2634_));
 sky130_fd_sc_hd__nand3_1 _6804_ (.A(_2469_),
    .B(_2470_),
    .C(_2634_),
    .Y(_2635_));
 sky130_fd_sc_hd__a21o_1 _6805_ (.A1(_2469_),
    .A2(_2470_),
    .B1(_2634_),
    .X(_2636_));
 sky130_fd_sc_hd__a21oi_1 _6806_ (.A1(_2635_),
    .A2(_2636_),
    .B1(_2473_),
    .Y(_2637_));
 sky130_fd_sc_hd__and3_1 _6807_ (.A(_2636_),
    .B(_2467_),
    .C(_2635_),
    .X(_2638_));
 sky130_fd_sc_hd__nand2_1 _6808_ (.A(_2558_),
    .B(_2562_),
    .Y(_2639_));
 sky130_fd_sc_hd__nand4_2 _6809_ (.A(_3021_),
    .B(net292),
    .C(net188),
    .D(net181),
    .Y(_2640_));
 sky130_fd_sc_hd__o2bb2ai_4 _6810_ (.A1_N(net292),
    .A2_N(net188),
    .B1(net302),
    .B2(_1953_),
    .Y(_2641_));
 sky130_fd_sc_hd__o2bb2ai_1 _6811_ (.A1_N(_2640_),
    .A2_N(_2641_),
    .B1(_2929_),
    .B2(_1643_),
    .Y(_2643_));
 sky130_fd_sc_hd__nand3b_2 _6812_ (.A_N(net302),
    .B(net292),
    .C(net187),
    .Y(_2644_));
 sky130_fd_sc_hd__o2111ai_4 _6813_ (.A1(_1985_),
    .A2(_2644_),
    .B1(net278),
    .C1(net193),
    .D1(_2641_),
    .Y(_2645_));
 sky130_fd_sc_hd__nand3_2 _6814_ (.A(_2639_),
    .B(_2643_),
    .C(_2645_),
    .Y(_2646_));
 sky130_fd_sc_hd__inv_2 _6815_ (.A(_2559_),
    .Y(_2647_));
 sky130_fd_sc_hd__o21a_1 _6816_ (.A1(_3381_),
    .A2(_2199_),
    .B1(_2558_),
    .X(_2648_));
 sky130_fd_sc_hd__a2bb2oi_1 _6817_ (.A1_N(_2928_),
    .A2_N(_1643_),
    .B1(_2640_),
    .B2(_2641_),
    .Y(_2649_));
 sky130_fd_sc_hd__and2_1 _6818_ (.A(net278),
    .B(net193),
    .X(_2650_));
 sky130_fd_sc_hd__and3_1 _6819_ (.A(_2641_),
    .B(_2650_),
    .C(_2640_),
    .X(_2651_));
 sky130_fd_sc_hd__o22ai_4 _6820_ (.A1(_2647_),
    .A2(_2648_),
    .B1(_2649_),
    .B2(_2651_),
    .Y(_2652_));
 sky130_fd_sc_hd__nand3_1 _6821_ (.A(net266),
    .B(net203),
    .C(net197),
    .Y(_2654_));
 sky130_fd_sc_hd__o21a_2 _6822_ (.A1(net203),
    .A2(net197),
    .B1(net266),
    .X(_2655_));
 sky130_fd_sc_hd__and3_1 _6823_ (.A(_2584_),
    .B(_2654_),
    .C(_2655_),
    .X(_2656_));
 sky130_fd_sc_hd__and3_2 _6824_ (.A(net268),
    .B(net203),
    .C(net197),
    .X(_2657_));
 sky130_fd_sc_hd__o21ai_4 _6825_ (.A1(net204),
    .A2(net197),
    .B1(net266),
    .Y(_2658_));
 sky130_fd_sc_hd__o22a_1 _6826_ (.A1(_3176_),
    .A2(_1394_),
    .B1(_2657_),
    .B2(_2658_),
    .X(_2659_));
 sky130_fd_sc_hd__o2bb2ai_2 _6827_ (.A1_N(_2646_),
    .A2_N(_2652_),
    .B1(_2656_),
    .B2(_2659_),
    .Y(_2660_));
 sky130_fd_sc_hd__nand4_2 _6828_ (.A(_2655_),
    .B(net212),
    .C(net266),
    .D(_2654_),
    .Y(_2661_));
 sky130_fd_sc_hd__o22ai_4 _6829_ (.A1(_3342_),
    .A2(_1394_),
    .B1(_2657_),
    .B2(_2658_),
    .Y(_2662_));
 sky130_fd_sc_hd__nand4_2 _6830_ (.A(_2646_),
    .B(_2652_),
    .C(_2661_),
    .D(_2662_),
    .Y(_2663_));
 sky130_fd_sc_hd__o21ai_1 _6831_ (.A1(_2575_),
    .A2(_2567_),
    .B1(_2580_),
    .Y(_2665_));
 sky130_fd_sc_hd__a21oi_1 _6832_ (.A1(_2660_),
    .A2(_2663_),
    .B1(_2665_),
    .Y(_2666_));
 sky130_fd_sc_hd__nand2_1 _6833_ (.A(_2560_),
    .B(_2562_),
    .Y(_2667_));
 sky130_fd_sc_hd__o22a_1 _6834_ (.A1(_1985_),
    .A2(_2478_),
    .B1(_2563_),
    .B2(_2564_),
    .X(_2668_));
 sky130_fd_sc_hd__a21oi_2 _6835_ (.A1(_2667_),
    .A2(_2668_),
    .B1(_2575_),
    .Y(_2669_));
 sky130_fd_sc_hd__o211a_1 _6836_ (.A1(_2568_),
    .A2(_2669_),
    .B1(_2663_),
    .C1(_2660_),
    .X(_2670_));
 sky130_fd_sc_hd__o22ai_2 _6837_ (.A1(_2637_),
    .A2(_2638_),
    .B1(_2666_),
    .B2(_2670_),
    .Y(_2671_));
 sky130_fd_sc_hd__inv_2 _6838_ (.A(_2663_),
    .Y(_2672_));
 sky130_fd_sc_hd__o21ai_4 _6839_ (.A1(_2568_),
    .A2(_2669_),
    .B1(_2660_),
    .Y(_2673_));
 sky130_fd_sc_hd__nor2_1 _6840_ (.A(_2637_),
    .B(_2638_),
    .Y(_2674_));
 sky130_fd_sc_hd__a21o_1 _6841_ (.A1(_2660_),
    .A2(_2663_),
    .B1(_2665_),
    .X(_2676_));
 sky130_fd_sc_hd__o211ai_4 _6842_ (.A1(_2672_),
    .A2(_2673_),
    .B1(_2674_),
    .C1(_2676_),
    .Y(_2677_));
 sky130_fd_sc_hd__nand2_1 _6843_ (.A(_2485_),
    .B(_2505_),
    .Y(_2678_));
 sky130_fd_sc_hd__nand2_1 _6844_ (.A(_2579_),
    .B(_2580_),
    .Y(_2679_));
 sky130_fd_sc_hd__a22oi_2 _6845_ (.A1(_2481_),
    .A2(_2678_),
    .B1(_2679_),
    .B2(_2587_),
    .Y(_2680_));
 sky130_fd_sc_hd__a22oi_2 _6846_ (.A1(_2680_),
    .A2(_2586_),
    .B1(_2582_),
    .B2(_2605_),
    .Y(_2681_));
 sky130_fd_sc_hd__a21oi_1 _6847_ (.A1(_2671_),
    .A2(_2677_),
    .B1(_2681_),
    .Y(_2682_));
 sky130_fd_sc_hd__and3_1 _6848_ (.A(_2671_),
    .B(_2677_),
    .C(_2681_),
    .X(_2683_));
 sky130_fd_sc_hd__o22ai_1 _6849_ (.A1(_2632_),
    .A2(_2633_),
    .B1(_2682_),
    .B2(_2683_),
    .Y(_2684_));
 sky130_fd_sc_hd__a21o_1 _6850_ (.A1(_2671_),
    .A2(_2677_),
    .B1(_2681_),
    .X(_2685_));
 sky130_fd_sc_hd__nand3_1 _6851_ (.A(_2671_),
    .B(_2677_),
    .C(_2681_),
    .Y(_2687_));
 sky130_fd_sc_hd__nor2_1 _6852_ (.A(_2632_),
    .B(_2633_),
    .Y(_2688_));
 sky130_fd_sc_hd__nand3_1 _6853_ (.A(_2685_),
    .B(_2687_),
    .C(_2688_),
    .Y(_2689_));
 sky130_fd_sc_hd__nand3b_2 _6854_ (.A_N(_2630_),
    .B(_2684_),
    .C(_2689_),
    .Y(_2690_));
 sky130_fd_sc_hd__o21ai_1 _6855_ (.A1(_2682_),
    .A2(_2683_),
    .B1(_2688_),
    .Y(_2691_));
 sky130_fd_sc_hd__o211ai_1 _6856_ (.A1(_2632_),
    .A2(_2633_),
    .B1(_2685_),
    .C1(_2687_),
    .Y(_2692_));
 sky130_fd_sc_hd__nand3_1 _6857_ (.A(_2691_),
    .B(_2630_),
    .C(_2692_),
    .Y(_2693_));
 sky130_fd_sc_hd__nand3_2 _6858_ (.A(_2690_),
    .B(_2613_),
    .C(_2693_),
    .Y(_2694_));
 sky130_fd_sc_hd__a21o_1 _6859_ (.A1(_2693_),
    .A2(_2690_),
    .B1(_2613_),
    .X(_2695_));
 sky130_fd_sc_hd__nand2_1 _6860_ (.A(_2618_),
    .B(_2624_),
    .Y(_2696_));
 sky130_fd_sc_hd__a21o_1 _6861_ (.A1(_2694_),
    .A2(_2695_),
    .B1(_2696_),
    .X(_2698_));
 sky130_fd_sc_hd__nand3_1 _6862_ (.A(_2696_),
    .B(_2695_),
    .C(_2694_),
    .Y(_2699_));
 sky130_fd_sc_hd__nand2_1 _6863_ (.A(_2698_),
    .B(_2699_),
    .Y(_2700_));
 sky130_fd_sc_hd__xnor2_1 _6864_ (.A(_2629_),
    .B(_2700_),
    .Y(_0096_));
 sky130_fd_sc_hd__a21oi_1 _6865_ (.A1(_2655_),
    .A2(net212),
    .B1(_2657_),
    .Y(_2701_));
 sky130_fd_sc_hd__o211ai_4 _6866_ (.A1(_2177_),
    .A2(_2382_),
    .B1(_2383_),
    .C1(_2701_),
    .Y(_2702_));
 sky130_fd_sc_hd__a31o_2 _6867_ (.A1(net266),
    .A2(net203),
    .A3(net198),
    .B1(net212),
    .X(_2703_));
 sky130_fd_sc_hd__nand4_4 _6868_ (.A(_2469_),
    .B(_2470_),
    .C(_2655_),
    .D(_2703_),
    .Y(_2704_));
 sky130_fd_sc_hd__and3_1 _6869_ (.A(_2702_),
    .B(_2704_),
    .C(_2473_),
    .X(_2705_));
 sky130_fd_sc_hd__a21oi_2 _6870_ (.A1(_2702_),
    .A2(_2704_),
    .B1(_2473_),
    .Y(_2706_));
 sky130_fd_sc_hd__nand4b_4 _6871_ (.A_N(net291),
    .B(net278),
    .C(net188),
    .D(net180),
    .Y(_2708_));
 sky130_fd_sc_hd__o2bb2ai_4 _6872_ (.A1_N(net278),
    .A2_N(net187),
    .B1(net291),
    .B2(_1958_),
    .Y(_2709_));
 sky130_fd_sc_hd__nand2_1 _6873_ (.A(net267),
    .B(net193),
    .Y(_2710_));
 sky130_fd_sc_hd__a21o_1 _6874_ (.A1(_2708_),
    .A2(_2709_),
    .B1(_2710_),
    .X(_2711_));
 sky130_fd_sc_hd__o211ai_2 _6875_ (.A1(_3058_),
    .A2(_1643_),
    .B1(_2708_),
    .C1(_2709_),
    .Y(_2712_));
 sky130_fd_sc_hd__a21boi_2 _6876_ (.A1(_2641_),
    .A2(_2650_),
    .B1_N(_2640_),
    .Y(_2713_));
 sky130_fd_sc_hd__and3_2 _6877_ (.A(_2711_),
    .B(_2712_),
    .C(_2713_),
    .X(_2714_));
 sky130_fd_sc_hd__o2bb2ai_2 _6878_ (.A1_N(_2650_),
    .A2_N(_2641_),
    .B1(_2644_),
    .B2(_1985_),
    .Y(_2715_));
 sky130_fd_sc_hd__o2bb2ai_2 _6879_ (.A1_N(_2708_),
    .A2_N(_2709_),
    .B1(_3058_),
    .B2(_1643_),
    .Y(_2716_));
 sky130_fd_sc_hd__nand4_2 _6880_ (.A(_2709_),
    .B(net193),
    .C(net267),
    .D(_2708_),
    .Y(_2717_));
 sky130_fd_sc_hd__nand3_2 _6881_ (.A(_2715_),
    .B(_2716_),
    .C(_2717_),
    .Y(_2719_));
 sky130_fd_sc_hd__o21ai_2 _6882_ (.A1(_2656_),
    .A2(_2659_),
    .B1(_2719_),
    .Y(_2720_));
 sky130_fd_sc_hd__o21ai_2 _6883_ (.A1(_2657_),
    .A2(_2658_),
    .B1(_2584_),
    .Y(_2721_));
 sky130_fd_sc_hd__o21ai_4 _6884_ (.A1(_2658_),
    .A2(_2703_),
    .B1(_2721_),
    .Y(_2722_));
 sky130_fd_sc_hd__a21boi_2 _6885_ (.A1(_2652_),
    .A2(_2722_),
    .B1_N(_2646_),
    .Y(_2723_));
 sky130_fd_sc_hd__nand3_1 _6886_ (.A(_1394_),
    .B(_2654_),
    .C(_2655_),
    .Y(_2724_));
 sky130_fd_sc_hd__nand3_2 _6887_ (.A(_2711_),
    .B(_2712_),
    .C(_2713_),
    .Y(_2725_));
 sky130_fd_sc_hd__a22o_1 _6888_ (.A1(_2721_),
    .A2(_2724_),
    .B1(_2725_),
    .B2(_2719_),
    .X(_2726_));
 sky130_fd_sc_hd__o211ai_4 _6889_ (.A1(_2714_),
    .A2(_2720_),
    .B1(_2723_),
    .C1(_2726_),
    .Y(_2727_));
 sky130_fd_sc_hd__nand2_2 _6890_ (.A(_2661_),
    .B(_2662_),
    .Y(_2728_));
 sky130_fd_sc_hd__a31o_1 _6891_ (.A1(_2715_),
    .A2(_2716_),
    .A3(_2717_),
    .B1(_2728_),
    .X(_2730_));
 sky130_fd_sc_hd__a22o_1 _6892_ (.A1(_2661_),
    .A2(_2662_),
    .B1(_2725_),
    .B2(_2719_),
    .X(_2731_));
 sky130_fd_sc_hd__a21oi_1 _6893_ (.A1(_2643_),
    .A2(_2645_),
    .B1(_2639_),
    .Y(_2732_));
 sky130_fd_sc_hd__o21ai_1 _6894_ (.A1(_2732_),
    .A2(_2728_),
    .B1(_2646_),
    .Y(_2733_));
 sky130_fd_sc_hd__o211ai_4 _6895_ (.A1(_2714_),
    .A2(_2730_),
    .B1(_2731_),
    .C1(_2733_),
    .Y(_2734_));
 sky130_fd_sc_hd__o211ai_2 _6896_ (.A1(_2705_),
    .A2(_2706_),
    .B1(_2727_),
    .C1(_2734_),
    .Y(_2735_));
 sky130_fd_sc_hd__nand3_1 _6897_ (.A(_2704_),
    .B(_2473_),
    .C(_2702_),
    .Y(_2736_));
 sky130_fd_sc_hd__a21o_1 _6898_ (.A1(_2702_),
    .A2(_2704_),
    .B1(_2473_),
    .X(_2737_));
 sky130_fd_sc_hd__nand2_2 _6899_ (.A(_2736_),
    .B(_2737_),
    .Y(_2738_));
 sky130_fd_sc_hd__a21o_1 _6900_ (.A1(_2727_),
    .A2(_2734_),
    .B1(_2738_),
    .X(_2739_));
 sky130_fd_sc_hd__o2111ai_4 _6901_ (.A1(_2673_),
    .A2(_2672_),
    .B1(_2735_),
    .C1(_2677_),
    .D1(_2739_),
    .Y(_2741_));
 sky130_fd_sc_hd__a21o_1 _6902_ (.A1(_2676_),
    .A2(_2674_),
    .B1(_2670_),
    .X(_2742_));
 sky130_fd_sc_hd__nor2_1 _6903_ (.A(_2705_),
    .B(_2706_),
    .Y(_2743_));
 sky130_fd_sc_hd__a21o_1 _6904_ (.A1(_2727_),
    .A2(_2734_),
    .B1(_2743_),
    .X(_2744_));
 sky130_fd_sc_hd__a31oi_2 _6905_ (.A1(_2715_),
    .A2(_2716_),
    .A3(_2717_),
    .B1(_2722_),
    .Y(_2745_));
 sky130_fd_sc_hd__nand2_1 _6906_ (.A(_2745_),
    .B(_2725_),
    .Y(_2746_));
 sky130_fd_sc_hd__a31oi_2 _6907_ (.A1(_2726_),
    .A2(_2723_),
    .A3(_2746_),
    .B1(_2738_),
    .Y(_2747_));
 sky130_fd_sc_hd__nand2_1 _6908_ (.A(_2747_),
    .B(_2734_),
    .Y(_2748_));
 sky130_fd_sc_hd__nand3_2 _6909_ (.A(_2742_),
    .B(_2744_),
    .C(_2748_),
    .Y(_2749_));
 sky130_fd_sc_hd__a31o_1 _6910_ (.A1(_2469_),
    .A2(_2470_),
    .A3(_2634_),
    .B1(_2638_),
    .X(_2750_));
 sky130_fd_sc_hd__xor2_2 _6911_ (.A(_2524_),
    .B(_2750_),
    .X(_2752_));
 sky130_fd_sc_hd__a21oi_1 _6912_ (.A1(_2741_),
    .A2(_2749_),
    .B1(_2752_),
    .Y(_2753_));
 sky130_fd_sc_hd__and3_1 _6913_ (.A(_2741_),
    .B(_2749_),
    .C(_2752_),
    .X(_2754_));
 sky130_fd_sc_hd__a21oi_1 _6914_ (.A1(_2685_),
    .A2(_2688_),
    .B1(_2683_),
    .Y(_2755_));
 sky130_fd_sc_hd__o21bai_1 _6915_ (.A1(_2753_),
    .A2(_2754_),
    .B1_N(_2755_),
    .Y(_2756_));
 sky130_fd_sc_hd__a21o_1 _6916_ (.A1(_2741_),
    .A2(_2749_),
    .B1(_2752_),
    .X(_2757_));
 sky130_fd_sc_hd__nand3_1 _6917_ (.A(_2741_),
    .B(_2749_),
    .C(_2752_),
    .Y(_2758_));
 sky130_fd_sc_hd__nand3_1 _6918_ (.A(_2757_),
    .B(_2758_),
    .C(_2755_),
    .Y(_2759_));
 sky130_fd_sc_hd__nand2_1 _6919_ (.A(_2756_),
    .B(_2759_),
    .Y(_2760_));
 sky130_fd_sc_hd__or2_1 _6920_ (.A(_2633_),
    .B(_2760_),
    .X(_2761_));
 sky130_fd_sc_hd__nand2_1 _6921_ (.A(_2760_),
    .B(_2633_),
    .Y(_2763_));
 sky130_fd_sc_hd__a22oi_2 _6922_ (.A1(_2690_),
    .A2(_2694_),
    .B1(_2761_),
    .B2(_2763_),
    .Y(_2764_));
 sky130_fd_sc_hd__nand4_1 _6923_ (.A(_2690_),
    .B(_2694_),
    .C(_2761_),
    .D(_2763_),
    .Y(_2765_));
 sky130_fd_sc_hd__nor2b_1 _6924_ (.A(_2764_),
    .B_N(_2765_),
    .Y(_2766_));
 sky130_fd_sc_hd__nor2_1 _6925_ (.A(_2628_),
    .B(_2700_),
    .Y(_2767_));
 sky130_fd_sc_hd__nand3_1 _6926_ (.A(_2461_),
    .B(_2551_),
    .C(_2767_),
    .Y(_2768_));
 sky130_fd_sc_hd__a21oi_1 _6927_ (.A1(_2694_),
    .A2(_2695_),
    .B1(_2696_),
    .Y(_2769_));
 sky130_fd_sc_hd__a21o_1 _6928_ (.A1(_2627_),
    .A2(_2699_),
    .B1(_2769_),
    .X(_2770_));
 sky130_fd_sc_hd__o31a_1 _6929_ (.A1(_2552_),
    .A2(_2628_),
    .A3(_2700_),
    .B1(_2770_),
    .X(_2771_));
 sky130_fd_sc_hd__nand2_1 _6930_ (.A(_2768_),
    .B(_2771_),
    .Y(_2772_));
 sky130_fd_sc_hd__xor2_1 _6931_ (.A(_2766_),
    .B(_2772_),
    .X(_0097_));
 sky130_fd_sc_hd__a21boi_1 _6932_ (.A1(_2749_),
    .A2(_2752_),
    .B1_N(_2741_),
    .Y(_2774_));
 sky130_fd_sc_hd__nand2_1 _6933_ (.A(_2704_),
    .B(_2736_),
    .Y(_2775_));
 sky130_fd_sc_hd__xor2_2 _6934_ (.A(_2524_),
    .B(_2775_),
    .X(_2776_));
 sky130_fd_sc_hd__o21ai_2 _6935_ (.A1(net192),
    .A2(net187),
    .B1(net267),
    .Y(_2777_));
 sky130_fd_sc_hd__and2_1 _6936_ (.A(net192),
    .B(net188),
    .X(_2778_));
 sky130_fd_sc_hd__o22ai_4 _6937_ (.A1(net278),
    .A2(_1958_),
    .B1(_2777_),
    .B2(_2778_),
    .Y(_2779_));
 sky130_fd_sc_hd__o21a_1 _6938_ (.A1(net193),
    .A2(net187),
    .B1(net267),
    .X(_2780_));
 sky130_fd_sc_hd__and2b_1 _6939_ (.A_N(net278),
    .B(net180),
    .X(_2781_));
 sky130_fd_sc_hd__nand2_1 _6940_ (.A(net193),
    .B(net187),
    .Y(_2782_));
 sky130_fd_sc_hd__nand3_2 _6941_ (.A(_2780_),
    .B(_2781_),
    .C(_2782_),
    .Y(_2784_));
 sky130_fd_sc_hd__nand2_1 _6942_ (.A(_2779_),
    .B(_2784_),
    .Y(_2785_));
 sky130_fd_sc_hd__o21ai_2 _6943_ (.A1(_3342_),
    .A2(_2199_),
    .B1(_2708_),
    .Y(_2786_));
 sky130_fd_sc_hd__nand2_1 _6944_ (.A(_2709_),
    .B(_2786_),
    .Y(_2787_));
 sky130_fd_sc_hd__nand2_1 _6945_ (.A(_2785_),
    .B(_2787_),
    .Y(_2788_));
 sky130_fd_sc_hd__nand4_2 _6946_ (.A(_2709_),
    .B(_2786_),
    .C(_2779_),
    .D(_2784_),
    .Y(_2789_));
 sky130_fd_sc_hd__and3_1 _6947_ (.A(_2722_),
    .B(_2788_),
    .C(_2789_),
    .X(_2790_));
 sky130_fd_sc_hd__and4_1 _6948_ (.A(_0509_),
    .B(net278),
    .C(net187),
    .D(net181),
    .X(_2791_));
 sky130_fd_sc_hd__a22oi_2 _6949_ (.A1(net278),
    .A2(net187),
    .B1(_0509_),
    .B2(net181),
    .Y(_2792_));
 sky130_fd_sc_hd__nor2_1 _6950_ (.A(_2710_),
    .B(_2792_),
    .Y(_2793_));
 sky130_fd_sc_hd__o21ai_1 _6951_ (.A1(_2791_),
    .A2(_2793_),
    .B1(_2785_),
    .Y(_2795_));
 sky130_fd_sc_hd__o2111ai_1 _6952_ (.A1(_2710_),
    .A2(_2792_),
    .B1(_2779_),
    .C1(_2784_),
    .D1(_2708_),
    .Y(_2796_));
 sky130_fd_sc_hd__nand3_1 _6953_ (.A(_2795_),
    .B(_2728_),
    .C(_2796_),
    .Y(_2797_));
 sky130_fd_sc_hd__nand3_2 _6954_ (.A(_2725_),
    .B(_2720_),
    .C(_2797_),
    .Y(_2798_));
 sky130_fd_sc_hd__nand3_1 _6955_ (.A(_2722_),
    .B(_2788_),
    .C(_2789_),
    .Y(_2799_));
 sky130_fd_sc_hd__nand2_1 _6956_ (.A(_2799_),
    .B(_2797_),
    .Y(_2800_));
 sky130_fd_sc_hd__o21ai_2 _6957_ (.A1(_2714_),
    .A2(_2745_),
    .B1(_2800_),
    .Y(_2801_));
 sky130_fd_sc_hd__o21a_1 _6958_ (.A1(_2790_),
    .A2(_2798_),
    .B1(_2801_),
    .X(_2802_));
 sky130_fd_sc_hd__o211ai_1 _6959_ (.A1(_2790_),
    .A2(_2798_),
    .B1(_2801_),
    .C1(_2738_),
    .Y(_2803_));
 sky130_fd_sc_hd__a21oi_1 _6960_ (.A1(_2746_),
    .A2(_2726_),
    .B1(_2723_),
    .Y(_2804_));
 sky130_fd_sc_hd__a21oi_1 _6961_ (.A1(_2727_),
    .A2(_2743_),
    .B1(_2804_),
    .Y(_2806_));
 sky130_fd_sc_hd__o211ai_2 _6962_ (.A1(_2738_),
    .A2(_2802_),
    .B1(_2803_),
    .C1(_2806_),
    .Y(_2807_));
 sky130_fd_sc_hd__o21ai_1 _6963_ (.A1(_2790_),
    .A2(_2798_),
    .B1(_2801_),
    .Y(_2808_));
 sky130_fd_sc_hd__o21ai_1 _6964_ (.A1(_2705_),
    .A2(_2706_),
    .B1(_2808_),
    .Y(_2809_));
 sky130_fd_sc_hd__o211ai_1 _6965_ (.A1(_2790_),
    .A2(_2798_),
    .B1(_2801_),
    .C1(_2743_),
    .Y(_2810_));
 sky130_fd_sc_hd__o211ai_2 _6966_ (.A1(_2804_),
    .A2(_2747_),
    .B1(_2809_),
    .C1(_2810_),
    .Y(_2811_));
 sky130_fd_sc_hd__nand3b_1 _6967_ (.A_N(_2776_),
    .B(_2807_),
    .C(_2811_),
    .Y(_2812_));
 sky130_fd_sc_hd__a21bo_1 _6968_ (.A1(_2807_),
    .A2(_2811_),
    .B1_N(_2776_),
    .X(_2813_));
 sky130_fd_sc_hd__nand3_1 _6969_ (.A(_2774_),
    .B(_2812_),
    .C(_2813_),
    .Y(_2814_));
 sky130_fd_sc_hd__a21o_1 _6970_ (.A1(_2812_),
    .A2(_2813_),
    .B1(_2774_),
    .X(_2815_));
 sky130_fd_sc_hd__o311a_1 _6971_ (.A1(net251),
    .A2(net244),
    .A3(net236),
    .B1(net266),
    .C1(_2750_),
    .X(_2817_));
 sky130_fd_sc_hd__a21bo_1 _6972_ (.A1(_2814_),
    .A2(_2815_),
    .B1_N(_2817_),
    .X(_2818_));
 sky130_fd_sc_hd__nand3b_1 _6973_ (.A_N(_2817_),
    .B(_2814_),
    .C(_2815_),
    .Y(_2819_));
 sky130_fd_sc_hd__a21oi_1 _6974_ (.A1(_2757_),
    .A2(_2758_),
    .B1(_2755_),
    .Y(_2820_));
 sky130_fd_sc_hd__a21oi_1 _6975_ (.A1(_2633_),
    .A2(_2759_),
    .B1(_2820_),
    .Y(_2821_));
 sky130_fd_sc_hd__a21oi_1 _6976_ (.A1(_2818_),
    .A2(_2819_),
    .B1(_2821_),
    .Y(_2822_));
 sky130_fd_sc_hd__and3_1 _6977_ (.A(_2818_),
    .B(_2819_),
    .C(_2821_),
    .X(_2823_));
 sky130_fd_sc_hd__nor2_1 _6978_ (.A(_2822_),
    .B(_2823_),
    .Y(_2824_));
 sky130_fd_sc_hd__o21ai_1 _6979_ (.A1(_2764_),
    .A2(_2772_),
    .B1(_2765_),
    .Y(_2825_));
 sky130_fd_sc_hd__xnor2_1 _6980_ (.A(_2824_),
    .B(_2825_),
    .Y(_0098_));
 sky130_fd_sc_hd__o311a_2 _6981_ (.A1(net251),
    .A2(net244),
    .A3(net236),
    .B1(net266),
    .C1(_2775_),
    .X(_2827_));
 sky130_fd_sc_hd__a31o_1 _6982_ (.A1(_2722_),
    .A2(_2788_),
    .A3(_2789_),
    .B1(_2798_),
    .X(_2828_));
 sky130_fd_sc_hd__nand2_1 _6983_ (.A(_2743_),
    .B(_2801_),
    .Y(_2829_));
 sky130_fd_sc_hd__o21ai_1 _6984_ (.A1(net267),
    .A2(_1985_),
    .B1(_2777_),
    .Y(_2830_));
 sky130_fd_sc_hd__nand2_1 _6985_ (.A(_2784_),
    .B(_2830_),
    .Y(_2831_));
 sky130_fd_sc_hd__nand2_1 _6986_ (.A(_2728_),
    .B(_2831_),
    .Y(_2832_));
 sky130_fd_sc_hd__a21o_1 _6987_ (.A1(_2721_),
    .A2(_2724_),
    .B1(_2831_),
    .X(_2833_));
 sky130_fd_sc_hd__nand2_1 _6988_ (.A(_2832_),
    .B(_2833_),
    .Y(_2834_));
 sky130_fd_sc_hd__o211ai_2 _6989_ (.A1(_2785_),
    .A2(_2787_),
    .B1(_2799_),
    .C1(_2834_),
    .Y(_2835_));
 sky130_fd_sc_hd__a22oi_1 _6990_ (.A1(_2709_),
    .A2(_2786_),
    .B1(_2779_),
    .B2(_2784_),
    .Y(_2836_));
 sky130_fd_sc_hd__o21ai_1 _6991_ (.A1(_2728_),
    .A2(_2836_),
    .B1(_2789_),
    .Y(_2838_));
 sky130_fd_sc_hd__nand3_1 _6992_ (.A(_2832_),
    .B(_2833_),
    .C(_2838_),
    .Y(_2839_));
 sky130_fd_sc_hd__a21o_1 _6993_ (.A1(_2835_),
    .A2(_2839_),
    .B1(_2738_),
    .X(_2840_));
 sky130_fd_sc_hd__o211ai_1 _6994_ (.A1(_2705_),
    .A2(_2706_),
    .B1(_2835_),
    .C1(_2839_),
    .Y(_2841_));
 sky130_fd_sc_hd__a22o_1 _6995_ (.A1(_2828_),
    .A2(_2829_),
    .B1(_2840_),
    .B2(_2841_),
    .X(_2842_));
 sky130_fd_sc_hd__nand4_1 _6996_ (.A(_2828_),
    .B(_2829_),
    .C(_2840_),
    .D(_2841_),
    .Y(_2843_));
 sky130_fd_sc_hd__a21oi_1 _6997_ (.A1(_2842_),
    .A2(_2843_),
    .B1(_2776_),
    .Y(_2844_));
 sky130_fd_sc_hd__nand3_1 _6998_ (.A(_2776_),
    .B(_2842_),
    .C(_2843_),
    .Y(_2845_));
 sky130_fd_sc_hd__and2b_1 _6999_ (.A_N(_2844_),
    .B(_2845_),
    .X(_2846_));
 sky130_fd_sc_hd__inv_2 _7000_ (.A(_2807_),
    .Y(_2847_));
 sky130_fd_sc_hd__o21ai_1 _7001_ (.A1(_2776_),
    .A2(_2847_),
    .B1(_2811_),
    .Y(_2849_));
 sky130_fd_sc_hd__xnor2_1 _7002_ (.A(_2846_),
    .B(_2849_),
    .Y(_2850_));
 sky130_fd_sc_hd__xnor2_1 _7003_ (.A(net941),
    .B(_2850_),
    .Y(_2851_));
 sky130_fd_sc_hd__a21boi_2 _7004_ (.A1(_2815_),
    .A2(net908),
    .B1_N(_2814_),
    .Y(_2852_));
 sky130_fd_sc_hd__xnor2_1 _7005_ (.A(_2851_),
    .B(_2852_),
    .Y(_2853_));
 sky130_fd_sc_hd__nand2_1 _7006_ (.A(_2552_),
    .B(_2770_),
    .Y(_2854_));
 sky130_fd_sc_hd__nand4_1 _7007_ (.A(_2258_),
    .B(_2049_),
    .C(_2048_),
    .D(_2043_),
    .Y(_2855_));
 sky130_fd_sc_hd__nand4_1 _7008_ (.A(_2457_),
    .B(_2548_),
    .C(_2550_),
    .D(_2358_),
    .Y(_2856_));
 sky130_fd_sc_hd__a21oi_1 _7009_ (.A1(_2460_),
    .A2(_2855_),
    .B1(_2856_),
    .Y(_2857_));
 sky130_fd_sc_hd__o21ai_1 _7010_ (.A1(_2628_),
    .A2(_2700_),
    .B1(_2770_),
    .Y(_2858_));
 sky130_fd_sc_hd__and3b_1 _7011_ (.A_N(_2764_),
    .B(_2824_),
    .C(_2765_),
    .X(_2860_));
 sky130_fd_sc_hd__o211ai_1 _7012_ (.A1(_2854_),
    .A2(_2857_),
    .B1(_2858_),
    .C1(_2860_),
    .Y(_2861_));
 sky130_fd_sc_hd__o21bai_1 _7013_ (.A1(_2764_),
    .A2(_2822_),
    .B1_N(_2823_),
    .Y(_2862_));
 sky130_fd_sc_hd__and3_1 _7014_ (.A(_2853_),
    .B(_2861_),
    .C(_2862_),
    .X(_2863_));
 sky130_fd_sc_hd__a21oi_1 _7015_ (.A1(_2861_),
    .A2(_2862_),
    .B1(_2853_),
    .Y(_2864_));
 sky130_fd_sc_hd__nor2_1 _7016_ (.A(_2863_),
    .B(_2864_),
    .Y(_0099_));
 sky130_fd_sc_hd__nor2_1 _7017_ (.A(_2851_),
    .B(_2852_),
    .Y(_2865_));
 sky130_fd_sc_hd__or2b_1 _7018_ (.A(_2846_),
    .B_N(_2849_),
    .X(_2866_));
 sky130_fd_sc_hd__a21boi_1 _7019_ (.A1(_2827_),
    .A2(_2850_),
    .B1_N(_2866_),
    .Y(_2867_));
 sky130_fd_sc_hd__mux2_1 _7020_ (.A0(_2843_),
    .A1(_2842_),
    .S(_2776_),
    .X(_2868_));
 sky130_fd_sc_hd__mux2_1 _7021_ (.A0(_2835_),
    .A1(_2839_),
    .S(_2738_),
    .X(_2870_));
 sky130_fd_sc_hd__xnor2_1 _7022_ (.A(_2827_),
    .B(_2832_),
    .Y(_2871_));
 sky130_fd_sc_hd__xnor2_1 _7023_ (.A(_2870_),
    .B(_2871_),
    .Y(_2872_));
 sky130_fd_sc_hd__xor2_1 _7024_ (.A(_2868_),
    .B(_2872_),
    .X(_2873_));
 sky130_fd_sc_hd__xnor2_1 _7025_ (.A(_2867_),
    .B(_2873_),
    .Y(_2874_));
 sky130_fd_sc_hd__o21bai_1 _7026_ (.A1(net909),
    .A2(_2864_),
    .B1_N(_2874_),
    .Y(_2875_));
 sky130_fd_sc_hd__inv_2 _7027_ (.A(_2862_),
    .Y(_2876_));
 sky130_fd_sc_hd__nand2_1 _7028_ (.A(_2766_),
    .B(_2824_),
    .Y(_2877_));
 sky130_fd_sc_hd__a21oi_1 _7029_ (.A1(_2768_),
    .A2(_2771_),
    .B1(_2877_),
    .Y(_2878_));
 sky130_fd_sc_hd__o21bai_1 _7030_ (.A1(_2876_),
    .A2(_2878_),
    .B1_N(_2853_),
    .Y(_2879_));
 sky130_fd_sc_hd__o211ai_1 _7031_ (.A1(_2851_),
    .A2(_2852_),
    .B1(_2874_),
    .C1(_2879_),
    .Y(_2881_));
 sky130_fd_sc_hd__nand2_1 _7032_ (.A(net910),
    .B(_2881_),
    .Y(_0100_));
 sky130_fd_sc_hd__and2b_1 _7033_ (.A_N(_1454_),
    .B(_1455_),
    .X(_2882_));
 sky130_fd_sc_hd__xnor2_1 _7034_ (.A(_1361_),
    .B(_2882_),
    .Y(_0086_));
 sky130_fd_sc_hd__o22a_1 _7035_ (.A1(_3178_),
    .A2(_2982_),
    .B1(_3295_),
    .B2(_1329_),
    .X(_2883_));
 sky130_fd_sc_hd__nor2_1 _7036_ (.A(_0425_),
    .B(_2883_),
    .Y(_0058_));
 sky130_fd_sc_hd__xor2_1 _7037_ (.A(_0425_),
    .B(_0429_),
    .X(_0059_));
 sky130_fd_sc_hd__o21ai_1 _7038_ (.A1(_0430_),
    .A2(_0432_),
    .B1(_0431_),
    .Y(_2884_));
 sky130_fd_sc_hd__xnor2_1 _7039_ (.A(_0395_),
    .B(_2884_),
    .Y(_0060_));
 sky130_fd_sc_hd__a311o_1 _7040_ (.A1(net386),
    .A2(net149),
    .A3(_0395_),
    .B1(_0403_),
    .C1(_0423_),
    .X(_2885_));
 sky130_fd_sc_hd__a21oi_1 _7041_ (.A1(_0435_),
    .A2(_2885_),
    .B1(_0433_),
    .Y(_2887_));
 sky130_fd_sc_hd__a21oi_1 _7042_ (.A1(_0435_),
    .A2(_0434_),
    .B1(_2887_),
    .Y(_0061_));
 sky130_fd_sc_hd__and2_1 _7043_ (.A(_0440_),
    .B(_0441_),
    .X(_2888_));
 sky130_fd_sc_hd__a21oi_1 _7044_ (.A1(_0400_),
    .A2(_0441_),
    .B1(_0440_),
    .Y(_2889_));
 sky130_fd_sc_hd__a21oi_1 _7045_ (.A1(_2888_),
    .A2(_0400_),
    .B1(_2889_),
    .Y(_0082_));
 sky130_fd_sc_hd__and3_1 _7046_ (.A(_0446_),
    .B(_0442_),
    .C(_0400_),
    .X(_2890_));
 sky130_fd_sc_hd__nor2_1 _7047_ (.A(_0447_),
    .B(_2890_),
    .Y(_0083_));
 sky130_fd_sc_hd__a22o_1 _7048_ (.A1(_0330_),
    .A2(_0332_),
    .B1(_0376_),
    .B2(_0443_),
    .X(_2891_));
 sky130_fd_sc_hd__or2_1 _7049_ (.A(_0447_),
    .B(_0378_),
    .X(_2892_));
 sky130_fd_sc_hd__and3_1 _7050_ (.A(_2891_),
    .B(_0448_),
    .C(_2892_),
    .X(_2893_));
 sky130_fd_sc_hd__clkbuf_1 _7051_ (.A(_2893_),
    .X(_0084_));
 sky130_fd_sc_hd__o21ai_1 _7052_ (.A1(_0322_),
    .A2(_0331_),
    .B1(_0321_),
    .Y(_2895_));
 sky130_fd_sc_hd__and4_1 _7053_ (.A(_0329_),
    .B(_2895_),
    .C(_0325_),
    .D(_0326_),
    .X(_2896_));
 sky130_fd_sc_hd__a22o_1 _7054_ (.A1(_0329_),
    .A2(_2895_),
    .B1(_0325_),
    .B2(_0326_),
    .X(_2897_));
 sky130_fd_sc_hd__a21o_1 _7055_ (.A1(_2891_),
    .A2(_0448_),
    .B1(_2897_),
    .X(_2898_));
 sky130_fd_sc_hd__a32oi_2 _7056_ (.A1(_2896_),
    .A2(_2891_),
    .A3(_0448_),
    .B1(_2898_),
    .B2(_0452_),
    .Y(_0085_));
 sky130_fd_sc_hd__nand2_1 _7057_ (.A(_0257_),
    .B(_0264_),
    .Y(_2899_));
 sky130_fd_sc_hd__xnor2_1 _7058_ (.A(_0452_),
    .B(_2899_),
    .Y(_0068_));
 sky130_fd_sc_hd__a21bo_1 _7059_ (.A1(_0452_),
    .A2(_0257_),
    .B1_N(_0264_),
    .X(_2900_));
 sky130_fd_sc_hd__o21ai_1 _7060_ (.A1(_0186_),
    .A2(_0187_),
    .B1(_0259_),
    .Y(_2901_));
 sky130_fd_sc_hd__xnor2_1 _7061_ (.A(_2900_),
    .B(_2901_),
    .Y(_0069_));
 sky130_fd_sc_hd__nand2_1 _7062_ (.A(_3505_),
    .B(_3506_),
    .Y(_2903_));
 sky130_fd_sc_hd__xor2_1 _7063_ (.A(_0453_),
    .B(_2903_),
    .X(_0070_));
 sky130_fd_sc_hd__nand2_1 _7064_ (.A(_0116_),
    .B(_0119_),
    .Y(_2904_));
 sky130_fd_sc_hd__a21boi_1 _7065_ (.A1(_0453_),
    .A2(_3506_),
    .B1_N(_3505_),
    .Y(_2905_));
 sky130_fd_sc_hd__xnor2_1 _7066_ (.A(_2904_),
    .B(_2905_),
    .Y(_0071_));
 sky130_fd_sc_hd__o2bb2a_1 _7067_ (.A1_N(_0116_),
    .A2_N(_0454_),
    .B1(_0120_),
    .B2(_0453_),
    .X(_2906_));
 sky130_fd_sc_hd__and2b_1 _7068_ (.A_N(_0483_),
    .B(_0477_),
    .X(_2907_));
 sky130_fd_sc_hd__xnor2_1 _7069_ (.A(_2906_),
    .B(_2907_),
    .Y(_0072_));
 sky130_fd_sc_hd__or2b_1 _7070_ (.A(_0479_),
    .B_N(_0472_),
    .X(_2908_));
 sky130_fd_sc_hd__o21a_1 _7071_ (.A1(_0483_),
    .A2(_2906_),
    .B1(_0477_),
    .X(_2910_));
 sky130_fd_sc_hd__xor2_1 _7072_ (.A(_2908_),
    .B(_2910_),
    .X(_0073_));
 sky130_fd_sc_hd__nand2_1 _7073_ (.A(_0482_),
    .B(_0484_),
    .Y(_2911_));
 sky130_fd_sc_hd__xnor2_2 _7074_ (.A(_0488_),
    .B(_2911_),
    .Y(_0074_));
 sky130_fd_sc_hd__a32oi_4 _7075_ (.A1(_0482_),
    .A2(_0484_),
    .A3(_0488_),
    .B1(_3088_),
    .B2(_0493_),
    .Y(_2912_));
 sky130_fd_sc_hd__a21oi_4 _7076_ (.A1(_3181_),
    .A2(_2912_),
    .B1(_0495_),
    .Y(_0075_));
 sky130_fd_sc_hd__dfrtp_1 _7077_ (.CLK(clknet_leaf_59_clk),
    .D(net509),
    .RESET_B(net464),
    .Q(\mixer_i.nco_valid ));
 sky130_fd_sc_hd__dfrtp_1 _7078_ (.CLK(clknet_leaf_59_clk),
    .D(_0025_),
    .RESET_B(net464),
    .Q(\nco_inst.phase_accum[0] ));
 sky130_fd_sc_hd__dfrtp_1 _7079_ (.CLK(clknet_leaf_59_clk),
    .D(net536),
    .RESET_B(net464),
    .Q(\nco_inst.phase_accum[1] ));
 sky130_fd_sc_hd__dfrtp_1 _7080_ (.CLK(clknet_leaf_60_clk),
    .D(net548),
    .RESET_B(net464),
    .Q(\nco_inst.phase_accum[2] ));
 sky130_fd_sc_hd__dfrtp_1 _7081_ (.CLK(clknet_leaf_60_clk),
    .D(net540),
    .RESET_B(net464),
    .Q(\nco_inst.phase_accum[3] ));
 sky130_fd_sc_hd__dfrtp_1 _7082_ (.CLK(clknet_leaf_60_clk),
    .D(net573),
    .RESET_B(net464),
    .Q(\nco_inst.phase_accum[4] ));
 sky130_fd_sc_hd__dfrtp_1 _7083_ (.CLK(clknet_leaf_61_clk),
    .D(net562),
    .RESET_B(net464),
    .Q(\nco_inst.phase_accum[5] ));
 sky130_fd_sc_hd__dfrtp_1 _7084_ (.CLK(clknet_leaf_61_clk),
    .D(net558),
    .RESET_B(net465),
    .Q(\nco_inst.phase_accum[6] ));
 sky130_fd_sc_hd__dfrtp_1 _7085_ (.CLK(clknet_leaf_61_clk),
    .D(net676),
    .RESET_B(net465),
    .Q(\nco_inst.phase_accum[7] ));
 sky130_fd_sc_hd__dfrtp_1 _7086_ (.CLK(clknet_leaf_0_clk),
    .D(net565),
    .RESET_B(net465),
    .Q(\nco_inst.phase_accum[8] ));
 sky130_fd_sc_hd__dfrtp_1 _7087_ (.CLK(clknet_leaf_0_clk),
    .D(net636),
    .RESET_B(net465),
    .Q(\nco_inst.phase_accum[9] ));
 sky130_fd_sc_hd__dfrtp_1 _7088_ (.CLK(clknet_leaf_0_clk),
    .D(net726),
    .RESET_B(net465),
    .Q(\nco_inst.phase_accum[10] ));
 sky130_fd_sc_hd__dfrtp_1 _7089_ (.CLK(clknet_leaf_0_clk),
    .D(net579),
    .RESET_B(net465),
    .Q(\nco_inst.phase_accum[11] ));
 sky130_fd_sc_hd__dfrtp_1 _7090_ (.CLK(clknet_leaf_1_clk),
    .D(net730),
    .RESET_B(net465),
    .Q(\nco_inst.phase_accum[12] ));
 sky130_fd_sc_hd__dfrtp_1 _7091_ (.CLK(clknet_leaf_1_clk),
    .D(net697),
    .RESET_B(net471),
    .Q(\nco_inst.phase_accum[13] ));
 sky130_fd_sc_hd__dfrtp_1 _7092_ (.CLK(clknet_leaf_1_clk),
    .D(net737),
    .RESET_B(net471),
    .Q(\nco_inst.phase_accum[14] ));
 sky130_fd_sc_hd__dfrtp_1 _7093_ (.CLK(clknet_leaf_9_clk),
    .D(net595),
    .RESET_B(net473),
    .Q(\nco_inst.phase_accum[15] ));
 sky130_fd_sc_hd__dfrtp_1 _7094_ (.CLK(clknet_leaf_9_clk),
    .D(net709),
    .RESET_B(net473),
    .Q(\nco_inst.phase_accum[16] ));
 sky130_fd_sc_hd__dfrtp_1 _7095_ (.CLK(clknet_leaf_9_clk),
    .D(net569),
    .RESET_B(net473),
    .Q(\nco_inst.phase_accum[17] ));
 sky130_fd_sc_hd__dfrtp_1 _7096_ (.CLK(clknet_leaf_10_clk),
    .D(_0034_),
    .RESET_B(net473),
    .Q(\nco_inst.phase_accum[18] ));
 sky130_fd_sc_hd__dfrtp_1 _7097_ (.CLK(clknet_leaf_10_clk),
    .D(net690),
    .RESET_B(net473),
    .Q(\nco_inst.phase_accum[19] ));
 sky130_fd_sc_hd__dfrtp_1 _7098_ (.CLK(clknet_leaf_11_clk),
    .D(net681),
    .RESET_B(net472),
    .Q(\nco_inst.phase_accum[20] ));
 sky130_fd_sc_hd__dfrtp_1 _7099_ (.CLK(clknet_leaf_11_clk),
    .D(net554),
    .RESET_B(net472),
    .Q(\nco_inst.phase_accum[21] ));
 sky130_fd_sc_hd__dfrtp_1 _7100_ (.CLK(clknet_leaf_11_clk),
    .D(net746),
    .RESET_B(net472),
    .Q(\nco_inst.phase_accum[22] ));
 sky130_fd_sc_hd__dfrtp_1 _7101_ (.CLK(clknet_leaf_11_clk),
    .D(net543),
    .RESET_B(net472),
    .Q(\nco_inst.phase_accum[23] ));
 sky130_fd_sc_hd__dfrtp_1 _7102_ (.CLK(clknet_leaf_11_clk),
    .D(net721),
    .RESET_B(net472),
    .Q(\nco_inst.cosine_lut.addr[0] ));
 sky130_fd_sc_hd__dfrtp_1 _7103_ (.CLK(clknet_leaf_11_clk),
    .D(net575),
    .RESET_B(net472),
    .Q(\nco_inst.cosine_lut.addr[1] ));
 sky130_fd_sc_hd__dfrtp_1 _7104_ (.CLK(clknet_leaf_12_clk),
    .D(_0043_),
    .RESET_B(net472),
    .Q(\nco_inst.cosine_lut.addr[2] ));
 sky130_fd_sc_hd__dfrtp_1 _7105_ (.CLK(clknet_leaf_12_clk),
    .D(net629),
    .RESET_B(net472),
    .Q(\nco_inst.cosine_lut.addr[3] ));
 sky130_fd_sc_hd__dfrtp_1 _7106_ (.CLK(clknet_leaf_12_clk),
    .D(net551),
    .RESET_B(net473),
    .Q(\nco_inst.cosine_lut.addr[4] ));
 sky130_fd_sc_hd__dfrtp_4 _7107_ (.CLK(clknet_leaf_12_clk),
    .D(net742),
    .RESET_B(net474),
    .Q(\nco_inst.cosine_lut.addr[5] ));
 sky130_fd_sc_hd__dfrtp_1 _7108_ (.CLK(clknet_leaf_12_clk),
    .D(net715),
    .RESET_B(net474),
    .Q(\nco_inst.lut_addr_sin[6] ));
 sky130_fd_sc_hd__dfrtp_1 _7109_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0049_),
    .RESET_B(net474),
    .Q(\nco_inst.lut_addr_sin[7] ));
 sky130_fd_sc_hd__dfrtp_1 _7110_ (.CLK(clknet_leaf_7_clk),
    .D(_0000_),
    .RESET_B(net478),
    .Q(\mixer_q.nco_data[0] ));
 sky130_fd_sc_hd__dfrtp_1 _7111_ (.CLK(clknet_leaf_8_clk),
    .D(_0003_),
    .RESET_B(net479),
    .Q(\mixer_q.nco_data[1] ));
 sky130_fd_sc_hd__dfrtp_1 _7112_ (.CLK(clknet_leaf_7_clk),
    .D(_0004_),
    .RESET_B(net478),
    .Q(\mixer_q.nco_data[2] ));
 sky130_fd_sc_hd__dfrtp_1 _7113_ (.CLK(clknet_leaf_8_clk),
    .D(_0005_),
    .RESET_B(net479),
    .Q(\mixer_q.nco_data[3] ));
 sky130_fd_sc_hd__dfrtp_1 _7114_ (.CLK(clknet_leaf_6_clk),
    .D(_0006_),
    .RESET_B(net476),
    .Q(\mixer_q.nco_data[4] ));
 sky130_fd_sc_hd__dfrtp_1 _7115_ (.CLK(clknet_leaf_2_clk),
    .D(_0007_),
    .RESET_B(net466),
    .Q(\mixer_q.nco_data[5] ));
 sky130_fd_sc_hd__dfrtp_1 _7116_ (.CLK(clknet_leaf_2_clk),
    .D(_0008_),
    .RESET_B(net466),
    .Q(\mixer_q.nco_data[6] ));
 sky130_fd_sc_hd__dfrtp_1 _7117_ (.CLK(clknet_leaf_2_clk),
    .D(_0009_),
    .RESET_B(net466),
    .Q(\mixer_q.nco_data[7] ));
 sky130_fd_sc_hd__dfrtp_1 _7118_ (.CLK(clknet_leaf_2_clk),
    .D(_0010_),
    .RESET_B(net466),
    .Q(\mixer_q.nco_data[8] ));
 sky130_fd_sc_hd__dfrtp_1 _7119_ (.CLK(clknet_leaf_2_clk),
    .D(_0011_),
    .RESET_B(net468),
    .Q(\mixer_q.nco_data[9] ));
 sky130_fd_sc_hd__dfrtp_1 _7120_ (.CLK(clknet_leaf_2_clk),
    .D(_0001_),
    .RESET_B(net466),
    .Q(\mixer_q.nco_data[10] ));
 sky130_fd_sc_hd__dfrtp_1 _7121_ (.CLK(clknet_leaf_2_clk),
    .D(_0002_),
    .RESET_B(net468),
    .Q(\mixer_q.nco_data[11] ));
 sky130_fd_sc_hd__dfrtp_4 _7122_ (.CLK(clknet_3_5__leaf_clk),
    .D(net177),
    .RESET_B(net486),
    .Q(\mixer_i.valid_stage2 ));
 sky130_fd_sc_hd__dfrtp_1 _7123_ (.CLK(clknet_leaf_50_clk),
    .D(_0062_),
    .RESET_B(net486),
    .Q(\mixer_i.product[0] ));
 sky130_fd_sc_hd__dfrtp_1 _7124_ (.CLK(clknet_leaf_45_clk),
    .D(_0063_),
    .RESET_B(net488),
    .Q(\mixer_i.product[1] ));
 sky130_fd_sc_hd__dfrtp_1 _7125_ (.CLK(clknet_leaf_48_clk),
    .D(_0064_),
    .RESET_B(net486),
    .Q(\mixer_i.product[2] ));
 sky130_fd_sc_hd__dfrtp_1 _7126_ (.CLK(clknet_leaf_48_clk),
    .D(_0065_),
    .RESET_B(net486),
    .Q(\mixer_i.product[3] ));
 sky130_fd_sc_hd__dfrtp_1 _7127_ (.CLK(clknet_leaf_46_clk),
    .D(_0066_),
    .RESET_B(net487),
    .Q(\mixer_i.product[4] ));
 sky130_fd_sc_hd__dfrtp_1 _7128_ (.CLK(clknet_leaf_45_clk),
    .D(_0086_),
    .RESET_B(net487),
    .Q(\mixer_i.product[5] ));
 sky130_fd_sc_hd__dfrtp_1 _7129_ (.CLK(clknet_leaf_46_clk),
    .D(_0101_),
    .RESET_B(net487),
    .Q(\mixer_i.product[6] ));
 sky130_fd_sc_hd__dfrtp_1 _7130_ (.CLK(clknet_leaf_42_clk),
    .D(_0102_),
    .RESET_B(net490),
    .Q(\mixer_i.product[7] ));
 sky130_fd_sc_hd__dfrtp_1 _7131_ (.CLK(clknet_leaf_42_clk),
    .D(_0103_),
    .RESET_B(net490),
    .Q(\mixer_i.product[8] ));
 sky130_fd_sc_hd__dfrtp_1 _7132_ (.CLK(clknet_leaf_42_clk),
    .D(_0104_),
    .RESET_B(net490),
    .Q(\mixer_i.product[9] ));
 sky130_fd_sc_hd__dfrtp_1 _7133_ (.CLK(clknet_leaf_41_clk),
    .D(_0087_),
    .RESET_B(net491),
    .Q(\mixer_i.product[10] ));
 sky130_fd_sc_hd__dfrtp_1 _7134_ (.CLK(clknet_leaf_41_clk),
    .D(_0088_),
    .RESET_B(net490),
    .Q(\mixer_i.product[11] ));
 sky130_fd_sc_hd__dfrtp_1 _7135_ (.CLK(clknet_leaf_39_clk),
    .D(_0089_),
    .RESET_B(net492),
    .Q(\mixer_i.product[12] ));
 sky130_fd_sc_hd__dfrtp_1 _7136_ (.CLK(clknet_leaf_39_clk),
    .D(_0090_),
    .RESET_B(net492),
    .Q(\mixer_i.product[13] ));
 sky130_fd_sc_hd__dfrtp_1 _7137_ (.CLK(clknet_leaf_35_clk),
    .D(_0091_),
    .RESET_B(net497),
    .Q(\mixer_i.product[14] ));
 sky130_fd_sc_hd__dfrtp_1 _7138_ (.CLK(clknet_leaf_35_clk),
    .D(_0092_),
    .RESET_B(net497),
    .Q(\mixer_i.product[15] ));
 sky130_fd_sc_hd__dfrtp_1 _7139_ (.CLK(clknet_leaf_33_clk),
    .D(_0093_),
    .RESET_B(net498),
    .Q(\mixer_i.product[16] ));
 sky130_fd_sc_hd__dfrtp_1 _7140_ (.CLK(clknet_leaf_34_clk),
    .D(_0094_),
    .RESET_B(net497),
    .Q(\mixer_i.product[17] ));
 sky130_fd_sc_hd__dfrtp_1 _7141_ (.CLK(clknet_leaf_33_clk),
    .D(_0095_),
    .RESET_B(net498),
    .Q(\mixer_i.product[18] ));
 sky130_fd_sc_hd__dfrtp_1 _7142_ (.CLK(clknet_leaf_33_clk),
    .D(_0096_),
    .RESET_B(net498),
    .Q(\mixer_i.product[19] ));
 sky130_fd_sc_hd__dfrtp_1 _7143_ (.CLK(clknet_leaf_31_clk),
    .D(_0097_),
    .RESET_B(net498),
    .Q(\mixer_i.product[20] ));
 sky130_fd_sc_hd__dfrtp_1 _7144_ (.CLK(clknet_leaf_31_clk),
    .D(_0098_),
    .RESET_B(net498),
    .Q(\mixer_i.product[21] ));
 sky130_fd_sc_hd__dfrtp_1 _7145_ (.CLK(clknet_leaf_31_clk),
    .D(_0099_),
    .RESET_B(net499),
    .Q(\mixer_i.product[22] ));
 sky130_fd_sc_hd__dfrtp_1 _7146_ (.CLK(clknet_leaf_31_clk),
    .D(net911),
    .RESET_B(net500),
    .Q(\mixer_i.product[23] ));
 sky130_fd_sc_hd__dfrtp_4 _7147_ (.CLK(clknet_leaf_58_clk),
    .D(net523),
    .RESET_B(net470),
    .Q(\mixer_i.adc_reg[0] ));
 sky130_fd_sc_hd__dfrtp_1 _7148_ (.CLK(clknet_leaf_58_clk),
    .D(net519),
    .RESET_B(net470),
    .Q(\mixer_i.adc_reg[1] ));
 sky130_fd_sc_hd__dfrtp_2 _7149_ (.CLK(clknet_leaf_57_clk),
    .D(net517),
    .RESET_B(net470),
    .Q(\mixer_i.adc_reg[2] ));
 sky130_fd_sc_hd__dfrtp_2 _7150_ (.CLK(clknet_leaf_57_clk),
    .D(net511),
    .RESET_B(net470),
    .Q(\mixer_i.adc_reg[3] ));
 sky130_fd_sc_hd__dfrtp_4 _7151_ (.CLK(clknet_leaf_57_clk),
    .D(net521),
    .RESET_B(net470),
    .Q(\mixer_i.adc_reg[4] ));
 sky130_fd_sc_hd__dfrtp_1 _7152_ (.CLK(clknet_leaf_57_clk),
    .D(net513),
    .RESET_B(net470),
    .Q(\mixer_i.adc_reg[5] ));
 sky130_fd_sc_hd__dfrtp_4 _7153_ (.CLK(clknet_3_4__leaf_clk),
    .D(net9),
    .RESET_B(net485),
    .Q(\mixer_i.adc_reg[6] ));
 sky130_fd_sc_hd__dfrtp_4 _7154_ (.CLK(clknet_3_4__leaf_clk),
    .D(net527),
    .RESET_B(net485),
    .Q(\mixer_i.adc_reg[7] ));
 sky130_fd_sc_hd__dfrtp_1 _7155_ (.CLK(clknet_3_4__leaf_clk),
    .D(net525),
    .RESET_B(net485),
    .Q(\mixer_i.adc_reg[8] ));
 sky130_fd_sc_hd__dfrtp_4 _7156_ (.CLK(clknet_3_4__leaf_clk),
    .D(net12),
    .RESET_B(net493),
    .Q(\mixer_i.adc_reg[9] ));
 sky130_fd_sc_hd__dfrtp_1 _7157_ (.CLK(clknet_3_5__leaf_clk),
    .D(net2),
    .RESET_B(net492),
    .Q(\mixer_i.adc_reg[10] ));
 sky130_fd_sc_hd__dfrtp_4 _7158_ (.CLK(clknet_leaf_40_clk),
    .D(net515),
    .RESET_B(net491),
    .Q(\mixer_i.adc_reg[11] ));
 sky130_fd_sc_hd__dfrtp_1 _7159_ (.CLK(clknet_leaf_28_clk),
    .D(net398),
    .RESET_B(net503),
    .Q(\mixer_i.valid_stage2_delayed ));
 sky130_fd_sc_hd__dfrtp_1 _7160_ (.CLK(clknet_3_6__leaf_clk),
    .D(net797),
    .RESET_B(net506),
    .Q(\mixer_i.nco_reg[0] ));
 sky130_fd_sc_hd__dfrtp_1 _7161_ (.CLK(clknet_3_6__leaf_clk),
    .D(net762),
    .RESET_B(net506),
    .Q(\mixer_i.nco_reg[1] ));
 sky130_fd_sc_hd__dfrtp_1 _7162_ (.CLK(clknet_3_6__leaf_clk),
    .D(net807),
    .RESET_B(net506),
    .Q(\mixer_i.nco_reg[2] ));
 sky130_fd_sc_hd__dfrtp_4 _7163_ (.CLK(clknet_leaf_7_clk),
    .D(net605),
    .RESET_B(net476),
    .Q(\mixer_i.nco_reg[3] ));
 sky130_fd_sc_hd__dfrtp_4 _7164_ (.CLK(clknet_leaf_5_clk),
    .D(net652),
    .RESET_B(net476),
    .Q(\mixer_i.nco_reg[4] ));
 sky130_fd_sc_hd__dfrtp_1 _7165_ (.CLK(clknet_leaf_38_clk),
    .D(net582),
    .RESET_B(net485),
    .Q(\mixer_i.nco_reg[5] ));
 sky130_fd_sc_hd__dfrtp_2 _7166_ (.CLK(clknet_leaf_55_clk),
    .D(net712),
    .RESET_B(net485),
    .Q(\mixer_i.nco_reg[6] ));
 sky130_fd_sc_hd__dfrtp_1 _7167_ (.CLK(clknet_leaf_38_clk),
    .D(net717),
    .RESET_B(net485),
    .Q(\mixer_i.nco_reg[7] ));
 sky130_fd_sc_hd__dfrtp_1 _7168_ (.CLK(clknet_leaf_55_clk),
    .D(net710),
    .RESET_B(net485),
    .Q(\mixer_i.nco_reg[8] ));
 sky130_fd_sc_hd__dfrtp_4 _7169_ (.CLK(clknet_leaf_3_clk),
    .D(net668),
    .RESET_B(net468),
    .Q(\mixer_i.nco_reg[9] ));
 sky130_fd_sc_hd__dfrtp_1 _7170_ (.CLK(clknet_leaf_38_clk),
    .D(net718),
    .RESET_B(net485),
    .Q(\mixer_i.nco_reg[10] ));
 sky130_fd_sc_hd__dfrtp_1 _7171_ (.CLK(clknet_leaf_38_clk),
    .D(net716),
    .RESET_B(net493),
    .Q(\mixer_i.nco_reg[11] ));
 sky130_fd_sc_hd__dfrtp_1 _7172_ (.CLK(clknet_leaf_50_clk),
    .D(net658),
    .RESET_B(net486),
    .Q(\mixer_i.product_delayed[0] ));
 sky130_fd_sc_hd__dfrtp_1 _7173_ (.CLK(clknet_leaf_47_clk),
    .D(net647),
    .RESET_B(net488),
    .Q(\mixer_i.product_delayed[1] ));
 sky130_fd_sc_hd__dfrtp_1 _7174_ (.CLK(clknet_leaf_49_clk),
    .D(net670),
    .RESET_B(net486),
    .Q(\mixer_i.product_delayed[2] ));
 sky130_fd_sc_hd__dfrtp_1 _7175_ (.CLK(clknet_leaf_48_clk),
    .D(net623),
    .RESET_B(net486),
    .Q(\mixer_i.product_delayed[3] ));
 sky130_fd_sc_hd__dfrtp_1 _7176_ (.CLK(clknet_leaf_46_clk),
    .D(net630),
    .RESET_B(net487),
    .Q(\mixer_i.product_delayed[4] ));
 sky130_fd_sc_hd__dfrtp_1 _7177_ (.CLK(clknet_leaf_46_clk),
    .D(net581),
    .RESET_B(net487),
    .Q(\mixer_i.product_delayed[5] ));
 sky130_fd_sc_hd__dfrtp_1 _7178_ (.CLK(clknet_leaf_46_clk),
    .D(net591),
    .RESET_B(net487),
    .Q(\mixer_i.product_delayed[6] ));
 sky130_fd_sc_hd__dfrtp_1 _7179_ (.CLK(clknet_leaf_42_clk),
    .D(net602),
    .RESET_B(net490),
    .Q(\mixer_i.product_delayed[7] ));
 sky130_fd_sc_hd__dfrtp_1 _7180_ (.CLK(clknet_leaf_42_clk),
    .D(net606),
    .RESET_B(net487),
    .Q(\mixer_i.product_delayed[8] ));
 sky130_fd_sc_hd__dfrtp_1 _7181_ (.CLK(clknet_leaf_40_clk),
    .D(net682),
    .RESET_B(net491),
    .Q(\mixer_i.product_delayed[9] ));
 sky130_fd_sc_hd__dfrtp_1 _7182_ (.CLK(clknet_leaf_41_clk),
    .D(net639),
    .RESET_B(net491),
    .Q(\mixer_i.product_delayed[10] ));
 sky130_fd_sc_hd__dfrtp_1 _7183_ (.CLK(clknet_leaf_41_clk),
    .D(net599),
    .RESET_B(net490),
    .Q(\mixer_i.product_delayed[11] ));
 sky130_fd_sc_hd__dfrtp_1 _7184_ (.CLK(clknet_leaf_39_clk),
    .D(net585),
    .RESET_B(net492),
    .Q(\mixer_i.product_delayed[12] ));
 sky130_fd_sc_hd__dfrtp_1 _7185_ (.CLK(clknet_leaf_35_clk),
    .D(net586),
    .RESET_B(net497),
    .Q(\mixer_i.product_delayed[13] ));
 sky130_fd_sc_hd__dfrtp_1 _7186_ (.CLK(clknet_leaf_35_clk),
    .D(net631),
    .RESET_B(net497),
    .Q(\mixer_i.product_delayed[14] ));
 sky130_fd_sc_hd__dfrtp_1 _7187_ (.CLK(clknet_leaf_35_clk),
    .D(net622),
    .RESET_B(net497),
    .Q(\mixer_i.product_delayed[15] ));
 sky130_fd_sc_hd__dfrtp_1 _7188_ (.CLK(clknet_leaf_32_clk),
    .D(net580),
    .RESET_B(net498),
    .Q(\mixer_i.product_delayed[16] ));
 sky130_fd_sc_hd__dfrtp_1 _7189_ (.CLK(clknet_leaf_34_clk),
    .D(net608),
    .RESET_B(net500),
    .Q(\mixer_i.product_delayed[17] ));
 sky130_fd_sc_hd__dfrtp_1 _7190_ (.CLK(clknet_leaf_32_clk),
    .D(net584),
    .RESET_B(net498),
    .Q(\mixer_i.product_delayed[18] ));
 sky130_fd_sc_hd__dfrtp_1 _7191_ (.CLK(clknet_leaf_30_clk),
    .D(net691),
    .RESET_B(net503),
    .Q(\mixer_i.product_delayed[19] ));
 sky130_fd_sc_hd__dfrtp_1 _7192_ (.CLK(clknet_leaf_29_clk),
    .D(net719),
    .RESET_B(net503),
    .Q(\mixer_i.product_delayed[20] ));
 sky130_fd_sc_hd__dfrtp_1 _7193_ (.CLK(clknet_leaf_29_clk),
    .D(net722),
    .RESET_B(net504),
    .Q(\mixer_i.product_delayed[21] ));
 sky130_fd_sc_hd__dfrtp_1 _7194_ (.CLK(clknet_leaf_30_clk),
    .D(net704),
    .RESET_B(net503),
    .Q(\mixer_i.product_delayed[22] ));
 sky130_fd_sc_hd__dfrtp_1 _7195_ (.CLK(clknet_leaf_31_clk),
    .D(net648),
    .RESET_B(net499),
    .Q(\mixer_i.product_delayed[23] ));
 sky130_fd_sc_hd__dfrtp_1 _7196_ (.CLK(clknet_leaf_50_clk),
    .D(net604),
    .RESET_B(net486),
    .Q(net47));
 sky130_fd_sc_hd__dfrtp_1 _7197_ (.CLK(clknet_leaf_50_clk),
    .D(net701),
    .RESET_B(net489),
    .Q(net58));
 sky130_fd_sc_hd__dfrtp_1 _7198_ (.CLK(clknet_leaf_49_clk),
    .D(net621),
    .RESET_B(net489),
    .Q(net63));
 sky130_fd_sc_hd__dfrtp_1 _7199_ (.CLK(clknet_leaf_48_clk),
    .D(net611),
    .RESET_B(net489),
    .Q(net64));
 sky130_fd_sc_hd__dfrtp_1 _7200_ (.CLK(clknet_leaf_47_clk),
    .D(net678),
    .RESET_B(net487),
    .Q(net65));
 sky130_fd_sc_hd__dfrtp_1 _7201_ (.CLK(clknet_leaf_46_clk),
    .D(net665),
    .RESET_B(net488),
    .Q(net66));
 sky130_fd_sc_hd__dfrtp_1 _7202_ (.CLK(clknet_leaf_46_clk),
    .D(net601),
    .RESET_B(net488),
    .Q(net67));
 sky130_fd_sc_hd__dfrtp_1 _7203_ (.CLK(clknet_leaf_42_clk),
    .D(net590),
    .RESET_B(net490),
    .Q(net68));
 sky130_fd_sc_hd__dfrtp_1 _7204_ (.CLK(clknet_leaf_42_clk),
    .D(net589),
    .RESET_B(net490),
    .Q(net69));
 sky130_fd_sc_hd__dfrtp_1 _7205_ (.CLK(clknet_leaf_40_clk),
    .D(net619),
    .RESET_B(net491),
    .Q(net70));
 sky130_fd_sc_hd__dfrtp_1 _7206_ (.CLK(clknet_leaf_40_clk),
    .D(net685),
    .RESET_B(net492),
    .Q(net48));
 sky130_fd_sc_hd__dfrtp_1 _7207_ (.CLK(clknet_leaf_41_clk),
    .D(net662),
    .RESET_B(net491),
    .Q(net49));
 sky130_fd_sc_hd__dfrtp_1 _7208_ (.CLK(clknet_leaf_39_clk),
    .D(net607),
    .RESET_B(net492),
    .Q(net50));
 sky130_fd_sc_hd__dfrtp_1 _7209_ (.CLK(clknet_leaf_35_clk),
    .D(net597),
    .RESET_B(net497),
    .Q(net51));
 sky130_fd_sc_hd__dfrtp_1 _7210_ (.CLK(clknet_leaf_34_clk),
    .D(net684),
    .RESET_B(net500),
    .Q(net52));
 sky130_fd_sc_hd__dfrtp_1 _7211_ (.CLK(clknet_leaf_35_clk),
    .D(net596),
    .RESET_B(net497),
    .Q(net53));
 sky130_fd_sc_hd__dfrtp_1 _7212_ (.CLK(clknet_leaf_32_clk),
    .D(net656),
    .RESET_B(net498),
    .Q(net54));
 sky130_fd_sc_hd__dfrtp_1 _7213_ (.CLK(clknet_leaf_32_clk),
    .D(net694),
    .RESET_B(net499),
    .Q(net55));
 sky130_fd_sc_hd__dfrtp_1 _7214_ (.CLK(clknet_leaf_30_clk),
    .D(net686),
    .RESET_B(net503),
    .Q(net56));
 sky130_fd_sc_hd__dfrtp_1 _7215_ (.CLK(clknet_leaf_30_clk),
    .D(net669),
    .RESET_B(net503),
    .Q(net57));
 sky130_fd_sc_hd__dfrtp_1 _7216_ (.CLK(clknet_leaf_29_clk),
    .D(net642),
    .RESET_B(net503),
    .Q(net59));
 sky130_fd_sc_hd__dfrtp_1 _7217_ (.CLK(clknet_leaf_29_clk),
    .D(net615),
    .RESET_B(net504),
    .Q(net60));
 sky130_fd_sc_hd__dfrtp_1 _7218_ (.CLK(clknet_leaf_30_clk),
    .D(net659),
    .RESET_B(net503),
    .Q(net61));
 sky130_fd_sc_hd__dfrtp_2 _7219_ (.CLK(clknet_leaf_31_clk),
    .D(net660),
    .RESET_B(net499),
    .Q(net62));
 sky130_fd_sc_hd__dfrtp_1 _7220_ (.CLK(clknet_leaf_28_clk),
    .D(net641),
    .RESET_B(net504),
    .Q(net95));
 sky130_fd_sc_hd__dfrtp_4 _7221_ (.CLK(clknet_leaf_59_clk),
    .D(_0024_),
    .RESET_B(net464),
    .Q(\mixer_i.valid_stage1 ));
 sky130_fd_sc_hd__dfrtp_1 _7222_ (.CLK(clknet_leaf_26_clk),
    .D(_0057_),
    .RESET_B(net501),
    .Q(\mixer_q.product[0] ));
 sky130_fd_sc_hd__dfrtp_1 _7223_ (.CLK(clknet_leaf_26_clk),
    .D(_0058_),
    .RESET_B(net501),
    .Q(\mixer_q.product[1] ));
 sky130_fd_sc_hd__dfrtp_1 _7224_ (.CLK(clknet_leaf_26_clk),
    .D(_0059_),
    .RESET_B(net501),
    .Q(\mixer_q.product[2] ));
 sky130_fd_sc_hd__dfrtp_1 _7225_ (.CLK(clknet_leaf_26_clk),
    .D(_0060_),
    .RESET_B(net501),
    .Q(\mixer_q.product[3] ));
 sky130_fd_sc_hd__dfrtp_1 _7226_ (.CLK(clknet_leaf_25_clk),
    .D(_0061_),
    .RESET_B(net494),
    .Q(\mixer_q.product[4] ));
 sky130_fd_sc_hd__dfrtp_1 _7227_ (.CLK(clknet_leaf_25_clk),
    .D(_0067_),
    .RESET_B(net494),
    .Q(\mixer_q.product[5] ));
 sky130_fd_sc_hd__dfrtp_1 _7228_ (.CLK(clknet_leaf_25_clk),
    .D(_0082_),
    .RESET_B(net495),
    .Q(\mixer_q.product[6] ));
 sky130_fd_sc_hd__dfrtp_1 _7229_ (.CLK(clknet_leaf_24_clk),
    .D(_0083_),
    .RESET_B(net494),
    .Q(\mixer_q.product[7] ));
 sky130_fd_sc_hd__dfrtp_1 _7230_ (.CLK(clknet_leaf_24_clk),
    .D(_0084_),
    .RESET_B(net494),
    .Q(\mixer_q.product[8] ));
 sky130_fd_sc_hd__dfrtp_1 _7231_ (.CLK(clknet_leaf_24_clk),
    .D(_0085_),
    .RESET_B(net494),
    .Q(\mixer_q.product[9] ));
 sky130_fd_sc_hd__dfrtp_1 _7232_ (.CLK(clknet_leaf_23_clk),
    .D(_0068_),
    .RESET_B(net496),
    .Q(\mixer_q.product[10] ));
 sky130_fd_sc_hd__dfrtp_1 _7233_ (.CLK(clknet_leaf_21_clk),
    .D(_0069_),
    .RESET_B(net482),
    .Q(\mixer_q.product[11] ));
 sky130_fd_sc_hd__dfrtp_1 _7234_ (.CLK(clknet_leaf_20_clk),
    .D(_0070_),
    .RESET_B(net482),
    .Q(\mixer_q.product[12] ));
 sky130_fd_sc_hd__dfrtp_1 _7235_ (.CLK(clknet_leaf_20_clk),
    .D(_0071_),
    .RESET_B(net482),
    .Q(\mixer_q.product[13] ));
 sky130_fd_sc_hd__dfrtp_1 _7236_ (.CLK(clknet_leaf_20_clk),
    .D(_0072_),
    .RESET_B(net480),
    .Q(\mixer_q.product[14] ));
 sky130_fd_sc_hd__dfrtp_1 _7237_ (.CLK(clknet_leaf_20_clk),
    .D(_0073_),
    .RESET_B(net480),
    .Q(\mixer_q.product[15] ));
 sky130_fd_sc_hd__dfrtp_1 _7238_ (.CLK(clknet_leaf_19_clk),
    .D(_0074_),
    .RESET_B(net480),
    .Q(\mixer_q.product[16] ));
 sky130_fd_sc_hd__dfrtp_1 _7239_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0075_),
    .RESET_B(net475),
    .Q(\mixer_q.product[17] ));
 sky130_fd_sc_hd__dfrtp_1 _7240_ (.CLK(clknet_leaf_7_clk),
    .D(_0076_),
    .RESET_B(net477),
    .Q(\mixer_q.product[18] ));
 sky130_fd_sc_hd__dfrtp_4 _7241_ (.CLK(clknet_leaf_5_clk),
    .D(_0077_),
    .RESET_B(net477),
    .Q(\mixer_q.product[19] ));
 sky130_fd_sc_hd__dfrtp_4 _7242_ (.CLK(clknet_leaf_5_clk),
    .D(_0078_),
    .RESET_B(net476),
    .Q(\mixer_q.product[20] ));
 sky130_fd_sc_hd__dfrtp_4 _7243_ (.CLK(clknet_leaf_5_clk),
    .D(_0079_),
    .RESET_B(net476),
    .Q(\mixer_q.product[21] ));
 sky130_fd_sc_hd__dfrtp_4 _7244_ (.CLK(clknet_leaf_4_clk),
    .D(_0080_),
    .RESET_B(net467),
    .Q(\mixer_q.product[22] ));
 sky130_fd_sc_hd__dfrtp_4 _7245_ (.CLK(clknet_leaf_2_clk),
    .D(_0081_),
    .RESET_B(net467),
    .Q(\mixer_q.product[23] ));
 sky130_fd_sc_hd__dfrtp_1 _7246_ (.CLK(clknet_leaf_7_clk),
    .D(net598),
    .RESET_B(net477),
    .Q(\mixer_q.nco_reg[0] ));
 sky130_fd_sc_hd__dfrtp_2 _7247_ (.CLK(clknet_leaf_8_clk),
    .D(net587),
    .RESET_B(net479),
    .Q(\mixer_q.nco_reg[1] ));
 sky130_fd_sc_hd__dfrtp_4 _7248_ (.CLK(clknet_leaf_5_clk),
    .D(net583),
    .RESET_B(net477),
    .Q(\mixer_q.nco_reg[2] ));
 sky130_fd_sc_hd__dfrtp_4 _7249_ (.CLK(clknet_leaf_8_clk),
    .D(net588),
    .RESET_B(net479),
    .Q(\mixer_q.nco_reg[3] ));
 sky130_fd_sc_hd__dfrtp_4 _7250_ (.CLK(clknet_leaf_6_clk),
    .D(net643),
    .RESET_B(net476),
    .Q(\mixer_q.nco_reg[4] ));
 sky130_fd_sc_hd__dfrtp_1 _7251_ (.CLK(clknet_leaf_4_clk),
    .D(net917),
    .RESET_B(net469),
    .Q(\mixer_q.nco_reg[5] ));
 sky130_fd_sc_hd__dfrtp_1 _7252_ (.CLK(clknet_leaf_2_clk),
    .D(net663),
    .RESET_B(net466),
    .Q(\mixer_q.nco_reg[6] ));
 sky130_fd_sc_hd__dfrtp_1 _7253_ (.CLK(clknet_leaf_2_clk),
    .D(net657),
    .RESET_B(net467),
    .Q(\mixer_q.nco_reg[7] ));
 sky130_fd_sc_hd__dfrtp_4 _7254_ (.CLK(clknet_leaf_4_clk),
    .D(net919),
    .RESET_B(net469),
    .Q(\mixer_q.nco_reg[8] ));
 sky130_fd_sc_hd__dfrtp_1 _7255_ (.CLK(clknet_leaf_3_clk),
    .D(net677),
    .RESET_B(net468),
    .Q(\mixer_q.nco_reg[9] ));
 sky130_fd_sc_hd__dfrtp_1 _7256_ (.CLK(clknet_leaf_56_clk),
    .D(net906),
    .RESET_B(net469),
    .Q(\mixer_q.nco_reg[10] ));
 sky130_fd_sc_hd__dfrtp_4 _7257_ (.CLK(clknet_leaf_56_clk),
    .D(net703),
    .RESET_B(net469),
    .Q(\mixer_q.nco_reg[11] ));
 sky130_fd_sc_hd__dfrtp_1 _7258_ (.CLK(clknet_leaf_26_clk),
    .D(net671),
    .RESET_B(net501),
    .Q(\mixer_q.product_delayed[0] ));
 sky130_fd_sc_hd__dfrtp_1 _7259_ (.CLK(clknet_leaf_27_clk),
    .D(net711),
    .RESET_B(net502),
    .Q(\mixer_q.product_delayed[1] ));
 sky130_fd_sc_hd__dfrtp_1 _7260_ (.CLK(clknet_leaf_26_clk),
    .D(net646),
    .RESET_B(net502),
    .Q(\mixer_q.product_delayed[2] ));
 sky130_fd_sc_hd__dfrtp_1 _7261_ (.CLK(clknet_leaf_26_clk),
    .D(net654),
    .RESET_B(net501),
    .Q(\mixer_q.product_delayed[3] ));
 sky130_fd_sc_hd__dfrtp_1 _7262_ (.CLK(clknet_leaf_26_clk),
    .D(net592),
    .RESET_B(net501),
    .Q(\mixer_q.product_delayed[4] ));
 sky130_fd_sc_hd__dfrtp_1 _7263_ (.CLK(clknet_leaf_25_clk),
    .D(net638),
    .RESET_B(net495),
    .Q(\mixer_q.product_delayed[5] ));
 sky130_fd_sc_hd__dfrtp_1 _7264_ (.CLK(clknet_leaf_25_clk),
    .D(net632),
    .RESET_B(net495),
    .Q(\mixer_q.product_delayed[6] ));
 sky130_fd_sc_hd__dfrtp_1 _7265_ (.CLK(clknet_leaf_24_clk),
    .D(net664),
    .RESET_B(net494),
    .Q(\mixer_q.product_delayed[7] ));
 sky130_fd_sc_hd__dfrtp_1 _7266_ (.CLK(clknet_leaf_24_clk),
    .D(net640),
    .RESET_B(net496),
    .Q(\mixer_q.product_delayed[8] ));
 sky130_fd_sc_hd__dfrtp_1 _7267_ (.CLK(clknet_leaf_23_clk),
    .D(net702),
    .RESET_B(net496),
    .Q(\mixer_q.product_delayed[9] ));
 sky130_fd_sc_hd__dfrtp_1 _7268_ (.CLK(clknet_leaf_23_clk),
    .D(net625),
    .RESET_B(net496),
    .Q(\mixer_q.product_delayed[10] ));
 sky130_fd_sc_hd__dfrtp_1 _7269_ (.CLK(clknet_leaf_21_clk),
    .D(net612),
    .RESET_B(net482),
    .Q(\mixer_q.product_delayed[11] ));
 sky130_fd_sc_hd__dfrtp_1 _7270_ (.CLK(clknet_leaf_21_clk),
    .D(net666),
    .RESET_B(net482),
    .Q(\mixer_q.product_delayed[12] ));
 sky130_fd_sc_hd__dfrtp_1 _7271_ (.CLK(clknet_leaf_20_clk),
    .D(net610),
    .RESET_B(net482),
    .Q(\mixer_q.product_delayed[13] ));
 sky130_fd_sc_hd__dfrtp_1 _7272_ (.CLK(clknet_leaf_20_clk),
    .D(net644),
    .RESET_B(net480),
    .Q(\mixer_q.product_delayed[14] ));
 sky130_fd_sc_hd__dfrtp_1 _7273_ (.CLK(clknet_leaf_19_clk),
    .D(net624),
    .RESET_B(net480),
    .Q(\mixer_q.product_delayed[15] ));
 sky130_fd_sc_hd__dfrtp_1 _7274_ (.CLK(clknet_leaf_19_clk),
    .D(net618),
    .RESET_B(net480),
    .Q(\mixer_q.product_delayed[16] ));
 sky130_fd_sc_hd__dfrtp_1 _7275_ (.CLK(clknet_leaf_19_clk),
    .D(net544),
    .RESET_B(net475),
    .Q(\mixer_q.product_delayed[17] ));
 sky130_fd_sc_hd__dfrtp_1 _7276_ (.CLK(clknet_leaf_18_clk),
    .D(net732),
    .RESET_B(net483),
    .Q(\mixer_q.product_delayed[18] ));
 sky130_fd_sc_hd__dfrtp_1 _7277_ (.CLK(clknet_leaf_16_clk),
    .D(net734),
    .RESET_B(net475),
    .Q(\mixer_q.product_delayed[19] ));
 sky130_fd_sc_hd__dfrtp_1 _7278_ (.CLK(clknet_leaf_19_clk),
    .D(net733),
    .RESET_B(net481),
    .Q(\mixer_q.product_delayed[20] ));
 sky130_fd_sc_hd__dfrtp_1 _7279_ (.CLK(clknet_leaf_15_clk),
    .D(net738),
    .RESET_B(net474),
    .Q(\mixer_q.product_delayed[21] ));
 sky130_fd_sc_hd__dfrtp_1 _7280_ (.CLK(clknet_leaf_14_clk),
    .D(net176),
    .RESET_B(net474),
    .Q(\mixer_q.product_delayed[22] ));
 sky130_fd_sc_hd__dfrtp_1 _7281_ (.CLK(clknet_leaf_14_clk),
    .D(net175),
    .RESET_B(net474),
    .Q(\mixer_q.product_delayed[23] ));
 sky130_fd_sc_hd__dfrtp_1 _7282_ (.CLK(clknet_leaf_27_clk),
    .D(net692),
    .RESET_B(net502),
    .Q(net71));
 sky130_fd_sc_hd__dfrtp_1 _7283_ (.CLK(clknet_leaf_27_clk),
    .D(net653),
    .RESET_B(net504),
    .Q(net82));
 sky130_fd_sc_hd__dfrtp_1 _7284_ (.CLK(clknet_leaf_27_clk),
    .D(net700),
    .RESET_B(net502),
    .Q(net87));
 sky130_fd_sc_hd__dfrtp_1 _7285_ (.CLK(clknet_leaf_26_clk),
    .D(net650),
    .RESET_B(net502),
    .Q(net88));
 sky130_fd_sc_hd__dfrtp_1 _7286_ (.CLK(clknet_leaf_26_clk),
    .D(net661),
    .RESET_B(net501),
    .Q(net89));
 sky130_fd_sc_hd__dfrtp_1 _7287_ (.CLK(clknet_leaf_25_clk),
    .D(net609),
    .RESET_B(net495),
    .Q(net90));
 sky130_fd_sc_hd__dfrtp_1 _7288_ (.CLK(clknet_leaf_25_clk),
    .D(net620),
    .RESET_B(net495),
    .Q(net91));
 sky130_fd_sc_hd__dfrtp_1 _7289_ (.CLK(clknet_leaf_24_clk),
    .D(net617),
    .RESET_B(net494),
    .Q(net92));
 sky130_fd_sc_hd__dfrtp_1 _7290_ (.CLK(clknet_leaf_24_clk),
    .D(net655),
    .RESET_B(net494),
    .Q(net93));
 sky130_fd_sc_hd__dfrtp_1 _7291_ (.CLK(clknet_leaf_24_clk),
    .D(net576),
    .RESET_B(net496),
    .Q(net94));
 sky130_fd_sc_hd__dfrtp_1 _7292_ (.CLK(clknet_leaf_23_clk),
    .D(net603),
    .RESET_B(net496),
    .Q(net72));
 sky130_fd_sc_hd__dfrtp_1 _7293_ (.CLK(clknet_leaf_23_clk),
    .D(net627),
    .RESET_B(net482),
    .Q(net73));
 sky130_fd_sc_hd__dfrtp_1 _7294_ (.CLK(clknet_leaf_21_clk),
    .D(net651),
    .RESET_B(net483),
    .Q(net74));
 sky130_fd_sc_hd__dfrtp_1 _7295_ (.CLK(clknet_leaf_20_clk),
    .D(net649),
    .RESET_B(net482),
    .Q(net75));
 sky130_fd_sc_hd__dfrtp_1 _7296_ (.CLK(clknet_leaf_20_clk),
    .D(net645),
    .RESET_B(net481),
    .Q(net76));
 sky130_fd_sc_hd__dfrtp_1 _7297_ (.CLK(clknet_leaf_19_clk),
    .D(net626),
    .RESET_B(net481),
    .Q(net77));
 sky130_fd_sc_hd__dfrtp_1 _7298_ (.CLK(clknet_leaf_19_clk),
    .D(net614),
    .RESET_B(net480),
    .Q(net78));
 sky130_fd_sc_hd__dfrtp_1 _7299_ (.CLK(clknet_leaf_16_clk),
    .D(net672),
    .RESET_B(net480),
    .Q(net79));
 sky130_fd_sc_hd__dfrtp_1 _7300_ (.CLK(clknet_leaf_18_clk),
    .D(net683),
    .RESET_B(net475),
    .Q(net80));
 sky130_fd_sc_hd__dfrtp_1 _7301_ (.CLK(clknet_leaf_16_clk),
    .D(net616),
    .RESET_B(net475),
    .Q(net81));
 sky130_fd_sc_hd__dfrtp_2 _7302_ (.CLK(clknet_leaf_20_clk),
    .D(net667),
    .RESET_B(net481),
    .Q(net83));
 sky130_fd_sc_hd__dfrtp_1 _7303_ (.CLK(clknet_leaf_15_clk),
    .D(net613),
    .RESET_B(net474),
    .Q(net84));
 sky130_fd_sc_hd__dfrtp_1 _7304_ (.CLK(clknet_leaf_14_clk),
    .D(net600),
    .RESET_B(net474),
    .Q(net85));
 sky130_fd_sc_hd__dfrtp_1 _7305_ (.CLK(clknet_leaf_14_clk),
    .D(net637),
    .RESET_B(net475),
    .Q(net86));
 sky130_fd_sc_hd__dfrtp_4 _7306_ (.CLK(clknet_leaf_7_clk),
    .D(_0012_),
    .RESET_B(net477),
    .Q(\mixer_i.nco_data[0] ));
 sky130_fd_sc_hd__dfrtp_2 _7307_ (.CLK(clknet_leaf_8_clk),
    .D(_0015_),
    .RESET_B(net479),
    .Q(\mixer_i.nco_data[1] ));
 sky130_fd_sc_hd__dfrtp_4 _7308_ (.CLK(clknet_leaf_6_clk),
    .D(_0016_),
    .RESET_B(net476),
    .Q(\mixer_i.nco_data[2] ));
 sky130_fd_sc_hd__dfrtp_1 _7309_ (.CLK(clknet_leaf_7_clk),
    .D(_0017_),
    .RESET_B(net477),
    .Q(\mixer_i.nco_data[3] ));
 sky130_fd_sc_hd__dfrtp_1 _7310_ (.CLK(clknet_leaf_6_clk),
    .D(_0018_),
    .RESET_B(net476),
    .Q(\mixer_i.nco_data[4] ));
 sky130_fd_sc_hd__dfrtp_1 _7311_ (.CLK(clknet_leaf_38_clk),
    .D(_0019_),
    .RESET_B(net493),
    .Q(\mixer_i.nco_data[5] ));
 sky130_fd_sc_hd__dfrtp_1 _7312_ (.CLK(clknet_leaf_3_clk),
    .D(_0020_),
    .RESET_B(net468),
    .Q(\mixer_i.nco_data[6] ));
 sky130_fd_sc_hd__dfrtp_1 _7313_ (.CLK(clknet_leaf_2_clk),
    .D(_0021_),
    .RESET_B(net467),
    .Q(\mixer_i.nco_data[7] ));
 sky130_fd_sc_hd__dfrtp_1 _7314_ (.CLK(clknet_leaf_3_clk),
    .D(_0022_),
    .RESET_B(net468),
    .Q(\mixer_i.nco_data[8] ));
 sky130_fd_sc_hd__dfrtp_1 _7315_ (.CLK(clknet_leaf_3_clk),
    .D(_0023_),
    .RESET_B(net468),
    .Q(\mixer_i.nco_data[9] ));
 sky130_fd_sc_hd__dfrtp_1 _7316_ (.CLK(clknet_leaf_2_clk),
    .D(_0013_),
    .RESET_B(net466),
    .Q(\mixer_i.nco_data[10] ));
 sky130_fd_sc_hd__dfrtp_1 _7317_ (.CLK(clknet_leaf_2_clk),
    .D(_0014_),
    .RESET_B(net466),
    .Q(\mixer_i.nco_data[11] ));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_0_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_Right_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_Right_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_Right_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_Right_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_Right_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_Right_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_Right_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_Right_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_Right_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_Right_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_Right_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_Right_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_Right_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_Right_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_Right_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_Right_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_Right_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_Right_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_120_Right_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_Right_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_Right_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_Right_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_124_Right_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_125_Right_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_126_Right_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_127_Right_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_128_Right_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_129_Right_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_130_Right_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_131_Right_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_132_Right_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_133_Right_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_134_Right_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_135_Right_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_136_Right_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_137_Right_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_138_Right_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_139_Right_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_140_Right_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_141_Right_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_142_Right_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_143_Right_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_144_Right_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_145_Right_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_146_Right_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_147_Right_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_148_Right_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_149_Right_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_150_Right_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_151_Right_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_152_Right_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_153_Right_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_154_Right_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_155_Right_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_156_Right_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_157_Right_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_158_Right_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_159_Right_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_160_Right_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_161_Right_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_162_Right_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_163_Right_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_164_Right_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_165_Right_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_166_Right_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_167_Right_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_168_Right_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_169_Right_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_170_Right_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_171_Right_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_172_Right_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_173_Right_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_174_Right_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_175_Right_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_176_Right_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_177_Right_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_178_Right_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_179_Right_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_180_Right_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_181_Right_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_182_Right_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_183_Right_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_184_Right_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_185_Right_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_186_Right_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_187_Right_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_188_Right_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_189_Right_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_190_Right_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_191_Right_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_192_Right_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_193_Right_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_194_Right_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_195_Right_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_196_Right_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_197_Right_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_198_Right_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_199_Right_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_200_Right_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_201_Right_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_202_Right_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_203_Right_203 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_204_Right_204 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_205_Right_205 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_206_Right_206 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_207_Right_207 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_208_Right_208 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_209_Right_209 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_210_Right_210 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_211_Right_211 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_212_Right_212 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_213_Right_213 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_214_Right_214 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_215_Right_215 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_216_Right_216 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_217_Right_217 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_218_Right_218 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_219_Right_219 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_220_Right_220 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_221_Right_221 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_222_Right_222 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_223_Right_223 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_224_Right_224 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_225_Right_225 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_226_Right_226 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_227 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_228 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_229 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_230 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_231 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_232 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_233 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_234 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_235 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_236 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_237 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_238 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_239 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_240 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_241 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_242 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_243 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_244 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_245 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_246 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_247 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_248 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_249 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_250 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_251 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_252 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_253 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_254 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_255 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_256 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_257 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_258 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_259 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_260 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_261 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_262 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_263 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_264 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_265 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_266 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_267 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_268 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_269 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_270 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_271 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_272 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_273 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_274 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_275 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_276 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_277 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_278 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_279 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_280 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_281 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_282 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_283 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_284 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_285 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_286 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_287 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_288 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_289 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_290 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_291 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_292 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_293 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_294 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_295 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_296 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_297 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_298 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_299 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_300 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_301 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_302 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_303 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_304 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_305 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_306 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_307 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_308 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_309 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_310 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_311 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_312 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_313 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_314 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_315 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_316 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_317 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_318 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_319 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_320 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_321 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_322 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_323 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_324 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_325 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_326 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_327 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_328 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_Left_329 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_Left_330 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_Left_331 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_Left_332 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_Left_333 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_Left_334 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_Left_335 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_Left_336 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_Left_337 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_Left_338 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_Left_339 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_Left_340 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_Left_341 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_Left_342 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_Left_343 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_Left_344 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_Left_345 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_Left_346 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_120_Left_347 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_Left_348 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_Left_349 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_Left_350 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_124_Left_351 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_125_Left_352 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_126_Left_353 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_127_Left_354 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_128_Left_355 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_129_Left_356 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_130_Left_357 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_131_Left_358 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_132_Left_359 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_133_Left_360 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_134_Left_361 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_135_Left_362 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_136_Left_363 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_137_Left_364 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_138_Left_365 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_139_Left_366 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_140_Left_367 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_141_Left_368 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_142_Left_369 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_143_Left_370 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_144_Left_371 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_145_Left_372 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_146_Left_373 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_147_Left_374 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_148_Left_375 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_149_Left_376 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_150_Left_377 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_151_Left_378 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_152_Left_379 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_153_Left_380 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_154_Left_381 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_155_Left_382 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_156_Left_383 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_157_Left_384 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_158_Left_385 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_159_Left_386 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_160_Left_387 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_161_Left_388 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_162_Left_389 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_163_Left_390 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_164_Left_391 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_165_Left_392 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_166_Left_393 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_167_Left_394 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_168_Left_395 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_169_Left_396 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_170_Left_397 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_171_Left_398 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_172_Left_399 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_173_Left_400 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_174_Left_401 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_175_Left_402 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_176_Left_403 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_177_Left_404 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_178_Left_405 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_179_Left_406 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_180_Left_407 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_181_Left_408 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_182_Left_409 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_183_Left_410 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_184_Left_411 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_185_Left_412 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_186_Left_413 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_187_Left_414 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_188_Left_415 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_189_Left_416 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_190_Left_417 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_191_Left_418 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_192_Left_419 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_193_Left_420 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_194_Left_421 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_195_Left_422 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_196_Left_423 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_197_Left_424 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_198_Left_425 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_199_Left_426 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_200_Left_427 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_201_Left_428 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_202_Left_429 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_203_Left_430 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_204_Left_431 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_205_Left_432 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_206_Left_433 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_207_Left_434 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_208_Left_435 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_209_Left_436 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_210_Left_437 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_211_Left_438 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_212_Left_439 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_213_Left_440 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_214_Left_441 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_215_Left_442 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_216_Left_443 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_217_Left_444 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_218_Left_445 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_219_Left_446 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_220_Left_447 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_221_Left_448 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_222_Left_449 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_223_Left_450 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_224_Left_451 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_225_Left_452 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_226_Left_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_5013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_5037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_5061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_5085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_5109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_5133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_5157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_5181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_5205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_5229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_5253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_5277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_5301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_5325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5949 ();
 sky130_fd_sc_hd__buf_2 input1 (.A(net522),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(net533),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(net514),
    .X(net3));
 sky130_fd_sc_hd__buf_2 input4 (.A(net518),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(net516),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(net510),
    .X(net6));
 sky130_fd_sc_hd__dlymetal6s2s_1 input7 (.A(net520),
    .X(net7));
 sky130_fd_sc_hd__buf_1 input8 (.A(net512),
    .X(net8));
 sky130_fd_sc_hd__buf_1 input9 (.A(net529),
    .X(net9));
 sky130_fd_sc_hd__buf_1 input10 (.A(net526),
    .X(net10));
 sky130_fd_sc_hd__buf_1 input11 (.A(net524),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 input12 (.A(net528),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(net530),
    .X(net13));
 sky130_fd_sc_hd__buf_1 input14 (.A(net534),
    .X(net14));
 sky130_fd_sc_hd__buf_1 input15 (.A(net723),
    .X(net15));
 sky130_fd_sc_hd__buf_1 input16 (.A(net577),
    .X(net16));
 sky130_fd_sc_hd__buf_1 input17 (.A(net727),
    .X(net17));
 sky130_fd_sc_hd__buf_1 input18 (.A(net695),
    .X(net18));
 sky130_fd_sc_hd__dlymetal6s2s_1 input19 (.A(net593),
    .X(net19));
 sky130_fd_sc_hd__buf_1 input20 (.A(net705),
    .X(net20));
 sky130_fd_sc_hd__buf_1 input21 (.A(net566),
    .X(net21));
 sky130_fd_sc_hd__buf_1 input22 (.A(net775),
    .X(net22));
 sky130_fd_sc_hd__buf_1 input23 (.A(phase_increment[18]),
    .X(net23));
 sky130_fd_sc_hd__buf_1 input24 (.A(net687),
    .X(net24));
 sky130_fd_sc_hd__buf_1 input25 (.A(net545),
    .X(net25));
 sky130_fd_sc_hd__dlymetal6s2s_1 input26 (.A(net679),
    .X(net26));
 sky130_fd_sc_hd__buf_1 input27 (.A(net552),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(net541),
    .X(net28));
 sky130_fd_sc_hd__buf_1 input29 (.A(phase_increment[23]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(net720),
    .X(net30));
 sky130_fd_sc_hd__dlymetal6s2s_1 input31 (.A(net574),
    .X(net31));
 sky130_fd_sc_hd__buf_1 input32 (.A(net802),
    .X(net32));
 sky130_fd_sc_hd__dlymetal6s2s_1 input33 (.A(net628),
    .X(net33));
 sky130_fd_sc_hd__buf_1 input34 (.A(net549),
    .X(net34));
 sky130_fd_sc_hd__dlymetal6s2s_1 input35 (.A(net741),
    .X(net35));
 sky130_fd_sc_hd__buf_1 input36 (.A(net537),
    .X(net36));
 sky130_fd_sc_hd__dlymetal6s2s_1 input37 (.A(net713),
    .X(net37));
 sky130_fd_sc_hd__buf_1 input38 (.A(net794),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(net570),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(net559),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(net555),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(phase_increment[6]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(net673),
    .X(net43));
 sky130_fd_sc_hd__buf_1 input44 (.A(net563),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(net633),
    .X(net45));
 sky130_fd_sc_hd__buf_1 input46 (.A(rst_n),
    .X(net46));
 sky130_fd_sc_hd__buf_8 output47 (.A(net774),
    .X(mixer_i_out[0]));
 sky130_fd_sc_hd__buf_8 output48 (.A(net769),
    .X(mixer_i_out[10]));
 sky130_fd_sc_hd__buf_8 output49 (.A(net805),
    .X(mixer_i_out[11]));
 sky130_fd_sc_hd__buf_8 output50 (.A(net750),
    .X(mixer_i_out[12]));
 sky130_fd_sc_hd__buf_8 output51 (.A(net949),
    .X(mixer_i_out[13]));
 sky130_fd_sc_hd__buf_8 output52 (.A(net752),
    .X(mixer_i_out[14]));
 sky130_fd_sc_hd__buf_8 output53 (.A(net791),
    .X(mixer_i_out[15]));
 sky130_fd_sc_hd__buf_8 output54 (.A(net758),
    .X(mixer_i_out[16]));
 sky130_fd_sc_hd__buf_8 output55 (.A(net761),
    .X(mixer_i_out[17]));
 sky130_fd_sc_hd__buf_8 output56 (.A(net766),
    .X(mixer_i_out[18]));
 sky130_fd_sc_hd__buf_8 output57 (.A(net765),
    .X(mixer_i_out[19]));
 sky130_fd_sc_hd__buf_8 output58 (.A(net784),
    .X(mixer_i_out[1]));
 sky130_fd_sc_hd__buf_8 output59 (.A(net759),
    .X(mixer_i_out[20]));
 sky130_fd_sc_hd__buf_8 output60 (.A(net768),
    .X(mixer_i_out[21]));
 sky130_fd_sc_hd__buf_8 output61 (.A(net799),
    .X(mixer_i_out[22]));
 sky130_fd_sc_hd__buf_8 output62 (.A(net808),
    .X(mixer_i_out[23]));
 sky130_fd_sc_hd__buf_8 output63 (.A(net767),
    .X(mixer_i_out[2]));
 sky130_fd_sc_hd__buf_8 output64 (.A(net783),
    .X(mixer_i_out[3]));
 sky130_fd_sc_hd__buf_8 output65 (.A(net770),
    .X(mixer_i_out[4]));
 sky130_fd_sc_hd__buf_8 output66 (.A(net771),
    .X(mixer_i_out[5]));
 sky130_fd_sc_hd__buf_8 output67 (.A(net780),
    .X(mixer_i_out[6]));
 sky130_fd_sc_hd__buf_8 output68 (.A(net773),
    .X(mixer_i_out[7]));
 sky130_fd_sc_hd__buf_8 output69 (.A(net789),
    .X(mixer_i_out[8]));
 sky130_fd_sc_hd__buf_8 output70 (.A(net782),
    .X(mixer_i_out[9]));
 sky130_fd_sc_hd__buf_8 output71 (.A(net804),
    .X(mixer_q_out[0]));
 sky130_fd_sc_hd__buf_8 output72 (.A(net753),
    .X(mixer_q_out[10]));
 sky130_fd_sc_hd__buf_8 output73 (.A(net760),
    .X(mixer_q_out[11]));
 sky130_fd_sc_hd__buf_8 output74 (.A(net763),
    .X(mixer_q_out[12]));
 sky130_fd_sc_hd__buf_8 output75 (.A(net764),
    .X(mixer_q_out[13]));
 sky130_fd_sc_hd__buf_8 output76 (.A(net757),
    .X(mixer_q_out[14]));
 sky130_fd_sc_hd__buf_8 output77 (.A(net755),
    .X(mixer_q_out[15]));
 sky130_fd_sc_hd__buf_8 output78 (.A(net756),
    .X(mixer_q_out[16]));
 sky130_fd_sc_hd__buf_8 output79 (.A(net747),
    .X(mixer_q_out[17]));
 sky130_fd_sc_hd__buf_8 output80 (.A(net796),
    .X(mixer_q_out[18]));
 sky130_fd_sc_hd__buf_8 output81 (.A(net748),
    .X(mixer_q_out[19]));
 sky130_fd_sc_hd__buf_8 output82 (.A(net772),
    .X(mixer_q_out[1]));
 sky130_fd_sc_hd__buf_8 output83 (.A(net806),
    .X(mixer_q_out[20]));
 sky130_fd_sc_hd__buf_8 output84 (.A(net740),
    .X(mixer_q_out[21]));
 sky130_fd_sc_hd__buf_8 output85 (.A(net749),
    .X(mixer_q_out[22]));
 sky130_fd_sc_hd__buf_8 output86 (.A(net751),
    .X(mixer_q_out[23]));
 sky130_fd_sc_hd__buf_8 output87 (.A(net781),
    .X(mixer_q_out[2]));
 sky130_fd_sc_hd__buf_8 output88 (.A(net800),
    .X(mixer_q_out[3]));
 sky130_fd_sc_hd__buf_8 output89 (.A(net798),
    .X(mixer_q_out[4]));
 sky130_fd_sc_hd__buf_8 output90 (.A(net793),
    .X(mixer_q_out[5]));
 sky130_fd_sc_hd__buf_8 output91 (.A(net785),
    .X(mixer_q_out[6]));
 sky130_fd_sc_hd__buf_8 output92 (.A(net790),
    .X(mixer_q_out[7]));
 sky130_fd_sc_hd__buf_8 output93 (.A(net788),
    .X(mixer_q_out[8]));
 sky130_fd_sc_hd__buf_8 output94 (.A(net792),
    .X(mixer_q_out[9]));
 sky130_fd_sc_hd__buf_8 output95 (.A(net754),
    .X(mixer_valid));
 sky130_fd_sc_hd__clkbuf_8 max_length96 (.A(_1793_),
    .X(net96));
 sky130_fd_sc_hd__buf_2 fanout97 (.A(net98),
    .X(net97));
 sky130_fd_sc_hd__buf_2 fanout98 (.A(net99),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_2 fanout99 (.A(net100),
    .X(net99));
 sky130_fd_sc_hd__buf_4 fanout100 (.A(\mixer_q.nco_reg[11] ),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_8 fanout101 (.A(\mixer_q.nco_reg[11] ),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_2 fanout102 (.A(\mixer_q.nco_reg[11] ),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_4 fanout103 (.A(net105),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_4 fanout104 (.A(net105),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_2 fanout105 (.A(net109),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_8 fanout106 (.A(net107),
    .X(net106));
 sky130_fd_sc_hd__buf_4 fanout107 (.A(net109),
    .X(net107));
 sky130_fd_sc_hd__buf_4 fanout108 (.A(net109),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_4 fanout109 (.A(\mixer_q.nco_reg[10] ),
    .X(net109));
 sky130_fd_sc_hd__buf_2 fanout110 (.A(net112),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_2 fanout111 (.A(net112),
    .X(net111));
 sky130_fd_sc_hd__buf_4 fanout112 (.A(net115),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_4 fanout113 (.A(net115),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_4 fanout114 (.A(net115),
    .X(net114));
 sky130_fd_sc_hd__buf_2 fanout115 (.A(\mixer_q.nco_reg[9] ),
    .X(net115));
 sky130_fd_sc_hd__buf_2 fanout116 (.A(net118),
    .X(net116));
 sky130_fd_sc_hd__buf_1 fanout117 (.A(net118),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_2 fanout118 (.A(net119),
    .X(net118));
 sky130_fd_sc_hd__buf_4 fanout119 (.A(\mixer_q.nco_reg[8] ),
    .X(net119));
 sky130_fd_sc_hd__buf_4 fanout120 (.A(net121),
    .X(net120));
 sky130_fd_sc_hd__buf_4 fanout121 (.A(\mixer_q.nco_reg[8] ),
    .X(net121));
 sky130_fd_sc_hd__buf_2 fanout122 (.A(net124),
    .X(net122));
 sky130_fd_sc_hd__buf_1 fanout123 (.A(net124),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_2 fanout124 (.A(net125),
    .X(net124));
 sky130_fd_sc_hd__buf_4 fanout125 (.A(net128),
    .X(net125));
 sky130_fd_sc_hd__buf_4 fanout126 (.A(net127),
    .X(net126));
 sky130_fd_sc_hd__buf_4 fanout127 (.A(net128),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_4 fanout128 (.A(\mixer_q.nco_reg[7] ),
    .X(net128));
 sky130_fd_sc_hd__buf_2 fanout129 (.A(net130),
    .X(net129));
 sky130_fd_sc_hd__buf_1 fanout130 (.A(net136),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_4 fanout131 (.A(net136),
    .X(net131));
 sky130_fd_sc_hd__buf_1 fanout132 (.A(net136),
    .X(net132));
 sky130_fd_sc_hd__buf_4 fanout133 (.A(net136),
    .X(net133));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout134 (.A(net135),
    .X(net134));
 sky130_fd_sc_hd__buf_4 fanout135 (.A(net136),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_4 fanout136 (.A(\mixer_q.nco_reg[6] ),
    .X(net136));
 sky130_fd_sc_hd__buf_2 fanout137 (.A(net143),
    .X(net137));
 sky130_fd_sc_hd__buf_1 fanout138 (.A(net143),
    .X(net138));
 sky130_fd_sc_hd__buf_4 fanout139 (.A(net140),
    .X(net139));
 sky130_fd_sc_hd__buf_4 fanout140 (.A(net143),
    .X(net140));
 sky130_fd_sc_hd__buf_2 fanout141 (.A(net143),
    .X(net141));
 sky130_fd_sc_hd__buf_2 fanout142 (.A(net143),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_4 fanout143 (.A(\mixer_q.nco_reg[5] ),
    .X(net143));
 sky130_fd_sc_hd__buf_2 fanout144 (.A(net145),
    .X(net144));
 sky130_fd_sc_hd__buf_2 fanout145 (.A(\mixer_q.nco_reg[4] ),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_4 fanout146 (.A(net150),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_4 fanout147 (.A(net150),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_4 fanout148 (.A(net150),
    .X(net148));
 sky130_fd_sc_hd__buf_2 fanout149 (.A(net150),
    .X(net149));
 sky130_fd_sc_hd__buf_2 fanout150 (.A(\mixer_q.nco_reg[4] ),
    .X(net150));
 sky130_fd_sc_hd__buf_2 fanout151 (.A(\mixer_q.nco_reg[3] ),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_4 fanout152 (.A(\mixer_q.nco_reg[3] ),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_4 fanout153 (.A(net155),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_2 fanout154 (.A(net155),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_4 fanout155 (.A(\mixer_q.nco_reg[3] ),
    .X(net155));
 sky130_fd_sc_hd__buf_2 fanout156 (.A(net157),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_2 fanout157 (.A(net158),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_4 fanout158 (.A(\mixer_q.nco_reg[2] ),
    .X(net158));
 sky130_fd_sc_hd__buf_4 fanout159 (.A(net160),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_2 fanout160 (.A(net162),
    .X(net160));
 sky130_fd_sc_hd__buf_2 fanout161 (.A(net162),
    .X(net161));
 sky130_fd_sc_hd__buf_2 fanout162 (.A(\mixer_q.nco_reg[2] ),
    .X(net162));
 sky130_fd_sc_hd__buf_2 fanout163 (.A(net164),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_2 fanout164 (.A(net165),
    .X(net164));
 sky130_fd_sc_hd__buf_4 fanout165 (.A(\mixer_q.nco_reg[1] ),
    .X(net165));
 sky130_fd_sc_hd__clkbuf_4 fanout166 (.A(net168),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_4 fanout167 (.A(net168),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_4 fanout168 (.A(net169),
    .X(net168));
 sky130_fd_sc_hd__buf_2 fanout169 (.A(\mixer_q.nco_reg[1] ),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_4 fanout170 (.A(net174),
    .X(net170));
 sky130_fd_sc_hd__buf_2 fanout171 (.A(net172),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_2 fanout172 (.A(net174),
    .X(net172));
 sky130_fd_sc_hd__buf_4 fanout173 (.A(net904),
    .X(net173));
 sky130_fd_sc_hd__buf_4 fanout174 (.A(\mixer_q.nco_reg[0] ),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_2 wire175 (.A(net810),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_2 wire176 (.A(net809),
    .X(net176));
 sky130_fd_sc_hd__buf_4 wire177 (.A(net811),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_4 fanout178 (.A(net179),
    .X(net178));
 sky130_fd_sc_hd__buf_6 fanout179 (.A(net181),
    .X(net179));
 sky130_fd_sc_hd__buf_4 fanout180 (.A(net181),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_4 fanout181 (.A(\mixer_i.nco_reg[11] ),
    .X(net181));
 sky130_fd_sc_hd__buf_4 fanout182 (.A(net184),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_2 fanout183 (.A(net184),
    .X(net183));
 sky130_fd_sc_hd__buf_4 fanout184 (.A(net189),
    .X(net184));
 sky130_fd_sc_hd__buf_4 fanout185 (.A(net189),
    .X(net185));
 sky130_fd_sc_hd__buf_2 fanout186 (.A(net189),
    .X(net186));
 sky130_fd_sc_hd__clkbuf_4 fanout187 (.A(net188),
    .X(net187));
 sky130_fd_sc_hd__buf_2 fanout188 (.A(net189),
    .X(net188));
 sky130_fd_sc_hd__clkbuf_2 fanout189 (.A(\mixer_i.nco_reg[10] ),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_4 fanout190 (.A(net191),
    .X(net190));
 sky130_fd_sc_hd__buf_2 fanout191 (.A(\mixer_i.nco_reg[9] ),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_4 fanout192 (.A(net194),
    .X(net192));
 sky130_fd_sc_hd__buf_2 fanout193 (.A(net194),
    .X(net193));
 sky130_fd_sc_hd__buf_2 fanout194 (.A(\mixer_i.nco_reg[9] ),
    .X(net194));
 sky130_fd_sc_hd__buf_4 fanout195 (.A(net200),
    .X(net195));
 sky130_fd_sc_hd__clkbuf_4 fanout196 (.A(net200),
    .X(net196));
 sky130_fd_sc_hd__buf_2 fanout197 (.A(net198),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_2 fanout198 (.A(net199),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_2 fanout199 (.A(net200),
    .X(net199));
 sky130_fd_sc_hd__buf_4 fanout200 (.A(\mixer_i.nco_reg[8] ),
    .X(net200));
 sky130_fd_sc_hd__buf_4 fanout201 (.A(net202),
    .X(net201));
 sky130_fd_sc_hd__clkbuf_4 fanout202 (.A(\mixer_i.nco_reg[7] ),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_2 fanout203 (.A(net204),
    .X(net203));
 sky130_fd_sc_hd__buf_2 fanout204 (.A(net205),
    .X(net204));
 sky130_fd_sc_hd__clkbuf_2 fanout205 (.A(net207),
    .X(net205));
 sky130_fd_sc_hd__clkbuf_4 fanout206 (.A(net207),
    .X(net206));
 sky130_fd_sc_hd__buf_2 fanout207 (.A(\mixer_i.nco_reg[7] ),
    .X(net207));
 sky130_fd_sc_hd__buf_4 fanout208 (.A(\mixer_i.nco_reg[6] ),
    .X(net208));
 sky130_fd_sc_hd__clkbuf_4 fanout209 (.A(\mixer_i.nco_reg[6] ),
    .X(net209));
 sky130_fd_sc_hd__buf_2 fanout210 (.A(net213),
    .X(net210));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout211 (.A(net213),
    .X(net211));
 sky130_fd_sc_hd__buf_2 fanout212 (.A(net213),
    .X(net212));
 sky130_fd_sc_hd__clkbuf_2 fanout213 (.A(\mixer_i.nco_reg[6] ),
    .X(net213));
 sky130_fd_sc_hd__buf_4 fanout214 (.A(net215),
    .X(net214));
 sky130_fd_sc_hd__buf_4 fanout215 (.A(net219),
    .X(net215));
 sky130_fd_sc_hd__buf_2 fanout216 (.A(net217),
    .X(net216));
 sky130_fd_sc_hd__clkbuf_2 fanout217 (.A(net218),
    .X(net217));
 sky130_fd_sc_hd__clkbuf_4 fanout218 (.A(net219),
    .X(net218));
 sky130_fd_sc_hd__buf_2 fanout219 (.A(\mixer_i.nco_reg[5] ),
    .X(net219));
 sky130_fd_sc_hd__buf_4 fanout220 (.A(net221),
    .X(net220));
 sky130_fd_sc_hd__buf_4 fanout221 (.A(net225),
    .X(net221));
 sky130_fd_sc_hd__buf_2 fanout222 (.A(net223),
    .X(net222));
 sky130_fd_sc_hd__clkbuf_2 fanout223 (.A(net224),
    .X(net223));
 sky130_fd_sc_hd__clkbuf_2 fanout224 (.A(net225),
    .X(net224));
 sky130_fd_sc_hd__clkbuf_4 fanout225 (.A(\mixer_i.nco_reg[4] ),
    .X(net225));
 sky130_fd_sc_hd__clkbuf_4 fanout226 (.A(net228),
    .X(net226));
 sky130_fd_sc_hd__clkbuf_4 fanout227 (.A(net228),
    .X(net227));
 sky130_fd_sc_hd__clkbuf_2 fanout228 (.A(\mixer_i.nco_reg[3] ),
    .X(net228));
 sky130_fd_sc_hd__clkbuf_4 fanout229 (.A(\mixer_i.nco_reg[3] ),
    .X(net229));
 sky130_fd_sc_hd__clkbuf_2 fanout230 (.A(\mixer_i.nco_reg[3] ),
    .X(net230));
 sky130_fd_sc_hd__clkbuf_2 fanout231 (.A(net232),
    .X(net231));
 sky130_fd_sc_hd__clkbuf_4 fanout232 (.A(net233),
    .X(net232));
 sky130_fd_sc_hd__buf_2 fanout233 (.A(net236),
    .X(net233));
 sky130_fd_sc_hd__clkbuf_4 fanout234 (.A(net235),
    .X(net234));
 sky130_fd_sc_hd__clkbuf_4 fanout235 (.A(net236),
    .X(net235));
 sky130_fd_sc_hd__clkbuf_4 fanout236 (.A(net907),
    .X(net236));
 sky130_fd_sc_hd__clkbuf_2 fanout237 (.A(net238),
    .X(net237));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout238 (.A(net239),
    .X(net238));
 sky130_fd_sc_hd__clkbuf_2 fanout239 (.A(net240),
    .X(net239));
 sky130_fd_sc_hd__buf_2 fanout240 (.A(net243),
    .X(net240));
 sky130_fd_sc_hd__clkbuf_2 fanout241 (.A(net242),
    .X(net241));
 sky130_fd_sc_hd__buf_4 fanout242 (.A(net243),
    .X(net242));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout243 (.A(net244),
    .X(net243));
 sky130_fd_sc_hd__buf_2 fanout244 (.A(net940),
    .X(net244));
 sky130_fd_sc_hd__buf_2 fanout245 (.A(net246),
    .X(net245));
 sky130_fd_sc_hd__clkbuf_2 fanout246 (.A(net247),
    .X(net246));
 sky130_fd_sc_hd__clkbuf_2 fanout247 (.A(net250),
    .X(net247));
 sky130_fd_sc_hd__buf_2 fanout248 (.A(net250),
    .X(net248));
 sky130_fd_sc_hd__clkbuf_2 fanout249 (.A(net250),
    .X(net249));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout250 (.A(net251),
    .X(net250));
 sky130_fd_sc_hd__clkbuf_4 fanout251 (.A(\mixer_i.nco_reg[0] ),
    .X(net251));
 sky130_fd_sc_hd__buf_2 fanout252 (.A(net255),
    .X(net252));
 sky130_fd_sc_hd__buf_2 fanout253 (.A(net255),
    .X(net253));
 sky130_fd_sc_hd__clkbuf_2 fanout254 (.A(net255),
    .X(net254));
 sky130_fd_sc_hd__clkbuf_2 fanout255 (.A(net260),
    .X(net255));
 sky130_fd_sc_hd__buf_2 fanout256 (.A(net258),
    .X(net256));
 sky130_fd_sc_hd__buf_1 fanout257 (.A(net258),
    .X(net257));
 sky130_fd_sc_hd__buf_2 fanout258 (.A(net259),
    .X(net258));
 sky130_fd_sc_hd__buf_2 fanout259 (.A(net260),
    .X(net259));
 sky130_fd_sc_hd__buf_2 fanout260 (.A(\mixer_i.adc_reg[11] ),
    .X(net260));
 sky130_fd_sc_hd__clkbuf_2 fanout261 (.A(net265),
    .X(net261));
 sky130_fd_sc_hd__buf_2 fanout262 (.A(net263),
    .X(net262));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout263 (.A(net264),
    .X(net263));
 sky130_fd_sc_hd__buf_2 fanout264 (.A(net265),
    .X(net264));
 sky130_fd_sc_hd__buf_1 fanout265 (.A(net268),
    .X(net265));
 sky130_fd_sc_hd__buf_2 fanout266 (.A(net268),
    .X(net266));
 sky130_fd_sc_hd__clkbuf_4 fanout267 (.A(net268),
    .X(net267));
 sky130_fd_sc_hd__buf_2 fanout268 (.A(\mixer_i.adc_reg[11] ),
    .X(net268));
 sky130_fd_sc_hd__buf_2 fanout269 (.A(net273),
    .X(net269));
 sky130_fd_sc_hd__clkbuf_2 fanout270 (.A(net273),
    .X(net270));
 sky130_fd_sc_hd__buf_4 fanout271 (.A(net272),
    .X(net271));
 sky130_fd_sc_hd__clkbuf_4 fanout272 (.A(net273),
    .X(net272));
 sky130_fd_sc_hd__buf_2 fanout273 (.A(net280),
    .X(net273));
 sky130_fd_sc_hd__clkbuf_2 fanout274 (.A(net275),
    .X(net274));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout275 (.A(net277),
    .X(net275));
 sky130_fd_sc_hd__buf_2 fanout276 (.A(net277),
    .X(net276));
 sky130_fd_sc_hd__clkbuf_2 fanout277 (.A(net280),
    .X(net277));
 sky130_fd_sc_hd__buf_4 fanout278 (.A(net280),
    .X(net278));
 sky130_fd_sc_hd__buf_2 fanout279 (.A(net280),
    .X(net279));
 sky130_fd_sc_hd__clkbuf_4 fanout280 (.A(\mixer_i.adc_reg[10] ),
    .X(net280));
 sky130_fd_sc_hd__buf_2 fanout281 (.A(net286),
    .X(net281));
 sky130_fd_sc_hd__clkbuf_2 fanout282 (.A(net286),
    .X(net282));
 sky130_fd_sc_hd__clkbuf_4 fanout283 (.A(net285),
    .X(net283));
 sky130_fd_sc_hd__clkbuf_4 fanout284 (.A(net285),
    .X(net284));
 sky130_fd_sc_hd__buf_4 fanout285 (.A(net286),
    .X(net285));
 sky130_fd_sc_hd__clkbuf_2 fanout286 (.A(\mixer_i.adc_reg[9] ),
    .X(net286));
 sky130_fd_sc_hd__clkbuf_4 fanout287 (.A(net289),
    .X(net287));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout288 (.A(net289),
    .X(net288));
 sky130_fd_sc_hd__clkbuf_4 fanout289 (.A(net293),
    .X(net289));
 sky130_fd_sc_hd__buf_2 fanout290 (.A(net291),
    .X(net290));
 sky130_fd_sc_hd__buf_2 fanout291 (.A(net292),
    .X(net291));
 sky130_fd_sc_hd__buf_2 fanout292 (.A(net293),
    .X(net292));
 sky130_fd_sc_hd__clkbuf_2 fanout293 (.A(\mixer_i.adc_reg[9] ),
    .X(net293));
 sky130_fd_sc_hd__buf_2 fanout294 (.A(net305),
    .X(net294));
 sky130_fd_sc_hd__buf_2 fanout295 (.A(net305),
    .X(net295));
 sky130_fd_sc_hd__clkbuf_4 fanout296 (.A(net298),
    .X(net296));
 sky130_fd_sc_hd__clkbuf_4 fanout297 (.A(net298),
    .X(net297));
 sky130_fd_sc_hd__buf_4 fanout298 (.A(net305),
    .X(net298));
 sky130_fd_sc_hd__clkbuf_4 fanout299 (.A(net301),
    .X(net299));
 sky130_fd_sc_hd__buf_2 fanout300 (.A(net301),
    .X(net300));
 sky130_fd_sc_hd__clkbuf_4 fanout301 (.A(net305),
    .X(net301));
 sky130_fd_sc_hd__buf_4 fanout302 (.A(net304),
    .X(net302));
 sky130_fd_sc_hd__buf_2 fanout303 (.A(net304),
    .X(net303));
 sky130_fd_sc_hd__buf_4 fanout304 (.A(net305),
    .X(net304));
 sky130_fd_sc_hd__clkbuf_4 fanout305 (.A(\mixer_i.adc_reg[8] ),
    .X(net305));
 sky130_fd_sc_hd__buf_4 fanout306 (.A(net308),
    .X(net306));
 sky130_fd_sc_hd__buf_4 fanout307 (.A(net308),
    .X(net307));
 sky130_fd_sc_hd__clkbuf_4 fanout308 (.A(net309),
    .X(net308));
 sky130_fd_sc_hd__buf_4 fanout309 (.A(\mixer_i.adc_reg[7] ),
    .X(net309));
 sky130_fd_sc_hd__clkbuf_4 fanout310 (.A(net315),
    .X(net310));
 sky130_fd_sc_hd__clkbuf_2 fanout311 (.A(net312),
    .X(net311));
 sky130_fd_sc_hd__clkbuf_4 fanout312 (.A(net315),
    .X(net312));
 sky130_fd_sc_hd__clkbuf_4 fanout313 (.A(net314),
    .X(net313));
 sky130_fd_sc_hd__clkbuf_4 fanout314 (.A(net315),
    .X(net314));
 sky130_fd_sc_hd__clkbuf_4 fanout315 (.A(\mixer_i.adc_reg[7] ),
    .X(net315));
 sky130_fd_sc_hd__clkbuf_4 fanout316 (.A(net317),
    .X(net316));
 sky130_fd_sc_hd__clkbuf_4 fanout317 (.A(net319),
    .X(net317));
 sky130_fd_sc_hd__buf_4 fanout318 (.A(net319),
    .X(net318));
 sky130_fd_sc_hd__buf_2 fanout319 (.A(net320),
    .X(net319));
 sky130_fd_sc_hd__clkbuf_4 fanout320 (.A(\mixer_i.adc_reg[6] ),
    .X(net320));
 sky130_fd_sc_hd__buf_4 fanout321 (.A(net324),
    .X(net321));
 sky130_fd_sc_hd__clkbuf_4 fanout322 (.A(net323),
    .X(net322));
 sky130_fd_sc_hd__buf_4 fanout323 (.A(net324),
    .X(net323));
 sky130_fd_sc_hd__buf_2 fanout324 (.A(net327),
    .X(net324));
 sky130_fd_sc_hd__clkbuf_4 fanout325 (.A(net327),
    .X(net325));
 sky130_fd_sc_hd__buf_4 fanout326 (.A(net327),
    .X(net326));
 sky130_fd_sc_hd__buf_2 fanout327 (.A(\mixer_i.adc_reg[6] ),
    .X(net327));
 sky130_fd_sc_hd__buf_2 fanout328 (.A(net329),
    .X(net328));
 sky130_fd_sc_hd__buf_4 fanout329 (.A(net330),
    .X(net329));
 sky130_fd_sc_hd__buf_4 fanout330 (.A(net331),
    .X(net330));
 sky130_fd_sc_hd__clkbuf_4 fanout331 (.A(net339),
    .X(net331));
 sky130_fd_sc_hd__buf_4 fanout332 (.A(net334),
    .X(net332));
 sky130_fd_sc_hd__clkbuf_2 fanout333 (.A(net334),
    .X(net333));
 sky130_fd_sc_hd__buf_2 fanout334 (.A(net339),
    .X(net334));
 sky130_fd_sc_hd__buf_4 fanout335 (.A(net336),
    .X(net335));
 sky130_fd_sc_hd__buf_4 fanout336 (.A(net339),
    .X(net336));
 sky130_fd_sc_hd__buf_4 fanout337 (.A(net338),
    .X(net337));
 sky130_fd_sc_hd__buf_4 fanout338 (.A(net339),
    .X(net338));
 sky130_fd_sc_hd__buf_4 fanout339 (.A(\mixer_i.adc_reg[5] ),
    .X(net339));
 sky130_fd_sc_hd__clkbuf_4 fanout340 (.A(net342),
    .X(net340));
 sky130_fd_sc_hd__clkbuf_4 fanout341 (.A(net342),
    .X(net341));
 sky130_fd_sc_hd__buf_2 fanout342 (.A(net345),
    .X(net342));
 sky130_fd_sc_hd__buf_2 fanout343 (.A(net344),
    .X(net343));
 sky130_fd_sc_hd__clkbuf_4 fanout344 (.A(net345),
    .X(net344));
 sky130_fd_sc_hd__buf_2 fanout345 (.A(\mixer_i.adc_reg[4] ),
    .X(net345));
 sky130_fd_sc_hd__buf_4 fanout346 (.A(net347),
    .X(net346));
 sky130_fd_sc_hd__clkbuf_4 fanout347 (.A(net348),
    .X(net347));
 sky130_fd_sc_hd__buf_2 fanout348 (.A(net350),
    .X(net348));
 sky130_fd_sc_hd__buf_4 fanout349 (.A(net350),
    .X(net349));
 sky130_fd_sc_hd__clkbuf_2 fanout350 (.A(net351),
    .X(net350));
 sky130_fd_sc_hd__clkbuf_8 fanout351 (.A(net352),
    .X(net351));
 sky130_fd_sc_hd__buf_4 wire352 (.A(\mixer_i.adc_reg[4] ),
    .X(net352));
 sky130_fd_sc_hd__buf_4 fanout353 (.A(net354),
    .X(net353));
 sky130_fd_sc_hd__buf_4 fanout354 (.A(net365),
    .X(net354));
 sky130_fd_sc_hd__clkbuf_4 fanout355 (.A(net356),
    .X(net355));
 sky130_fd_sc_hd__clkbuf_4 fanout356 (.A(net357),
    .X(net356));
 sky130_fd_sc_hd__clkbuf_2 fanout357 (.A(net365),
    .X(net357));
 sky130_fd_sc_hd__clkbuf_8 fanout358 (.A(net359),
    .X(net358));
 sky130_fd_sc_hd__clkbuf_4 fanout359 (.A(net362),
    .X(net359));
 sky130_fd_sc_hd__buf_4 fanout360 (.A(net362),
    .X(net360));
 sky130_fd_sc_hd__buf_2 fanout361 (.A(net362),
    .X(net361));
 sky130_fd_sc_hd__buf_2 fanout362 (.A(net365),
    .X(net362));
 sky130_fd_sc_hd__clkbuf_4 fanout363 (.A(net364),
    .X(net363));
 sky130_fd_sc_hd__buf_4 fanout364 (.A(net365),
    .X(net364));
 sky130_fd_sc_hd__buf_2 fanout365 (.A(\mixer_i.adc_reg[3] ),
    .X(net365));
 sky130_fd_sc_hd__buf_4 fanout366 (.A(net377),
    .X(net366));
 sky130_fd_sc_hd__buf_2 fanout367 (.A(net368),
    .X(net367));
 sky130_fd_sc_hd__clkbuf_2 fanout368 (.A(net370),
    .X(net368));
 sky130_fd_sc_hd__buf_4 fanout369 (.A(net370),
    .X(net369));
 sky130_fd_sc_hd__clkbuf_8 fanout370 (.A(net377),
    .X(net370));
 sky130_fd_sc_hd__buf_4 fanout371 (.A(net372),
    .X(net371));
 sky130_fd_sc_hd__buf_4 fanout372 (.A(net377),
    .X(net372));
 sky130_fd_sc_hd__buf_4 fanout373 (.A(net374),
    .X(net373));
 sky130_fd_sc_hd__buf_2 fanout374 (.A(net377),
    .X(net374));
 sky130_fd_sc_hd__clkbuf_4 fanout375 (.A(net376),
    .X(net375));
 sky130_fd_sc_hd__clkbuf_4 fanout376 (.A(net377),
    .X(net376));
 sky130_fd_sc_hd__buf_4 fanout377 (.A(\mixer_i.adc_reg[2] ),
    .X(net377));
 sky130_fd_sc_hd__clkbuf_4 fanout378 (.A(net389),
    .X(net378));
 sky130_fd_sc_hd__clkbuf_2 fanout379 (.A(net380),
    .X(net379));
 sky130_fd_sc_hd__buf_2 fanout380 (.A(net381),
    .X(net380));
 sky130_fd_sc_hd__clkbuf_4 fanout381 (.A(net389),
    .X(net381));
 sky130_fd_sc_hd__buf_4 fanout382 (.A(net385),
    .X(net382));
 sky130_fd_sc_hd__clkbuf_4 fanout383 (.A(net384),
    .X(net383));
 sky130_fd_sc_hd__buf_4 fanout384 (.A(net385),
    .X(net384));
 sky130_fd_sc_hd__buf_2 fanout385 (.A(net388),
    .X(net385));
 sky130_fd_sc_hd__buf_2 fanout386 (.A(net388),
    .X(net386));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout387 (.A(net388),
    .X(net387));
 sky130_fd_sc_hd__clkbuf_4 fanout388 (.A(net389),
    .X(net388));
 sky130_fd_sc_hd__clkbuf_4 fanout389 (.A(\mixer_i.adc_reg[1] ),
    .X(net389));
 sky130_fd_sc_hd__buf_2 fanout390 (.A(net391),
    .X(net390));
 sky130_fd_sc_hd__clkbuf_4 fanout391 (.A(net392),
    .X(net391));
 sky130_fd_sc_hd__clkbuf_4 fanout392 (.A(\mixer_i.adc_reg[0] ),
    .X(net392));
 sky130_fd_sc_hd__buf_4 fanout393 (.A(net395),
    .X(net393));
 sky130_fd_sc_hd__clkbuf_4 fanout394 (.A(net395),
    .X(net394));
 sky130_fd_sc_hd__buf_2 fanout395 (.A(net397),
    .X(net395));
 sky130_fd_sc_hd__clkbuf_4 fanout396 (.A(net397),
    .X(net396));
 sky130_fd_sc_hd__buf_2 fanout397 (.A(\mixer_i.adc_reg[0] ),
    .X(net397));
 sky130_fd_sc_hd__clkbuf_2 wire398 (.A(net739),
    .X(net398));
 sky130_fd_sc_hd__clkbuf_2 fanout399 (.A(net400),
    .X(net399));
 sky130_fd_sc_hd__clkbuf_2 fanout400 (.A(net401),
    .X(net400));
 sky130_fd_sc_hd__clkbuf_4 fanout401 (.A(net786),
    .X(net401));
 sky130_fd_sc_hd__buf_2 fanout402 (.A(net403),
    .X(net402));
 sky130_fd_sc_hd__clkbuf_2 fanout403 (.A(net405),
    .X(net403));
 sky130_fd_sc_hd__buf_2 fanout404 (.A(net405),
    .X(net404));
 sky130_fd_sc_hd__clkbuf_2 fanout405 (.A(net406),
    .X(net405));
 sky130_fd_sc_hd__buf_4 fanout406 (.A(net801),
    .X(net406));
 sky130_fd_sc_hd__buf_4 fanout407 (.A(net411),
    .X(net407));
 sky130_fd_sc_hd__buf_2 fanout408 (.A(net411),
    .X(net408));
 sky130_fd_sc_hd__buf_2 fanout409 (.A(net410),
    .X(net409));
 sky130_fd_sc_hd__clkbuf_4 fanout410 (.A(net411),
    .X(net410));
 sky130_fd_sc_hd__clkbuf_2 fanout411 (.A(\nco_inst.cosine_lut.addr[5] ),
    .X(net411));
 sky130_fd_sc_hd__buf_2 fanout412 (.A(net413),
    .X(net412));
 sky130_fd_sc_hd__clkbuf_4 fanout413 (.A(\nco_inst.cosine_lut.addr[5] ),
    .X(net413));
 sky130_fd_sc_hd__buf_4 fanout414 (.A(net419),
    .X(net414));
 sky130_fd_sc_hd__clkbuf_4 fanout415 (.A(net418),
    .X(net415));
 sky130_fd_sc_hd__clkbuf_2 fanout416 (.A(net418),
    .X(net416));
 sky130_fd_sc_hd__clkbuf_2 fanout417 (.A(net418),
    .X(net417));
 sky130_fd_sc_hd__clkbuf_2 fanout418 (.A(net419),
    .X(net418));
 sky130_fd_sc_hd__clkbuf_2 fanout419 (.A(net424),
    .X(net419));
 sky130_fd_sc_hd__clkbuf_4 fanout420 (.A(net424),
    .X(net420));
 sky130_fd_sc_hd__clkbuf_2 fanout421 (.A(net424),
    .X(net421));
 sky130_fd_sc_hd__clkbuf_4 fanout422 (.A(net423),
    .X(net422));
 sky130_fd_sc_hd__buf_2 fanout423 (.A(net424),
    .X(net423));
 sky130_fd_sc_hd__buf_2 fanout424 (.A(\nco_inst.cosine_lut.addr[4] ),
    .X(net424));
 sky130_fd_sc_hd__clkbuf_4 fanout425 (.A(net427),
    .X(net425));
 sky130_fd_sc_hd__clkbuf_4 fanout426 (.A(net427),
    .X(net426));
 sky130_fd_sc_hd__clkbuf_4 fanout427 (.A(net441),
    .X(net427));
 sky130_fd_sc_hd__buf_2 fanout428 (.A(net432),
    .X(net428));
 sky130_fd_sc_hd__clkbuf_2 fanout429 (.A(net432),
    .X(net429));
 sky130_fd_sc_hd__buf_2 fanout430 (.A(net432),
    .X(net430));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout431 (.A(net432),
    .X(net431));
 sky130_fd_sc_hd__clkbuf_2 fanout432 (.A(net441),
    .X(net432));
 sky130_fd_sc_hd__buf_2 fanout433 (.A(net435),
    .X(net433));
 sky130_fd_sc_hd__buf_1 fanout434 (.A(net435),
    .X(net434));
 sky130_fd_sc_hd__buf_2 fanout435 (.A(net436),
    .X(net435));
 sky130_fd_sc_hd__clkbuf_4 fanout436 (.A(net441),
    .X(net436));
 sky130_fd_sc_hd__clkbuf_4 fanout437 (.A(net440),
    .X(net437));
 sky130_fd_sc_hd__buf_2 fanout438 (.A(net440),
    .X(net438));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout439 (.A(net440),
    .X(net439));
 sky130_fd_sc_hd__buf_2 fanout440 (.A(net441),
    .X(net440));
 sky130_fd_sc_hd__buf_2 fanout441 (.A(\nco_inst.cosine_lut.addr[3] ),
    .X(net441));
 sky130_fd_sc_hd__clkbuf_4 fanout442 (.A(net450),
    .X(net442));
 sky130_fd_sc_hd__clkbuf_2 fanout443 (.A(net450),
    .X(net443));
 sky130_fd_sc_hd__buf_2 fanout444 (.A(net445),
    .X(net444));
 sky130_fd_sc_hd__buf_2 fanout445 (.A(net450),
    .X(net445));
 sky130_fd_sc_hd__buf_4 fanout446 (.A(net449),
    .X(net446));
 sky130_fd_sc_hd__clkbuf_2 fanout447 (.A(net449),
    .X(net447));
 sky130_fd_sc_hd__buf_2 fanout448 (.A(net449),
    .X(net448));
 sky130_fd_sc_hd__buf_2 fanout449 (.A(net450),
    .X(net449));
 sky130_fd_sc_hd__clkbuf_2 fanout450 (.A(\nco_inst.cosine_lut.addr[2] ),
    .X(net450));
 sky130_fd_sc_hd__buf_2 fanout451 (.A(net452),
    .X(net451));
 sky130_fd_sc_hd__clkbuf_4 fanout452 (.A(net457),
    .X(net452));
 sky130_fd_sc_hd__clkbuf_4 fanout453 (.A(net454),
    .X(net453));
 sky130_fd_sc_hd__buf_2 fanout454 (.A(net456),
    .X(net454));
 sky130_fd_sc_hd__buf_2 fanout455 (.A(net456),
    .X(net455));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout456 (.A(net457),
    .X(net456));
 sky130_fd_sc_hd__buf_2 fanout457 (.A(net914),
    .X(net457));
 sky130_fd_sc_hd__clkbuf_4 fanout458 (.A(net459),
    .X(net458));
 sky130_fd_sc_hd__clkbuf_4 fanout459 (.A(net463),
    .X(net459));
 sky130_fd_sc_hd__buf_2 fanout460 (.A(net461),
    .X(net460));
 sky130_fd_sc_hd__clkbuf_4 fanout461 (.A(net463),
    .X(net461));
 sky130_fd_sc_hd__clkbuf_4 fanout462 (.A(net463),
    .X(net462));
 sky130_fd_sc_hd__buf_2 fanout463 (.A(\nco_inst.cosine_lut.addr[0] ),
    .X(net463));
 sky130_fd_sc_hd__clkbuf_4 fanout464 (.A(net465),
    .X(net464));
 sky130_fd_sc_hd__clkbuf_4 fanout465 (.A(net471),
    .X(net465));
 sky130_fd_sc_hd__buf_2 fanout466 (.A(net468),
    .X(net466));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout467 (.A(net469),
    .X(net467));
 sky130_fd_sc_hd__buf_2 fanout468 (.A(net469),
    .X(net468));
 sky130_fd_sc_hd__buf_2 fanout469 (.A(net470),
    .X(net469));
 sky130_fd_sc_hd__clkbuf_4 fanout470 (.A(net471),
    .X(net470));
 sky130_fd_sc_hd__buf_4 fanout471 (.A(net507),
    .X(net471));
 sky130_fd_sc_hd__buf_2 fanout472 (.A(net473),
    .X(net472));
 sky130_fd_sc_hd__buf_2 fanout473 (.A(net484),
    .X(net473));
 sky130_fd_sc_hd__clkbuf_4 fanout474 (.A(net475),
    .X(net474));
 sky130_fd_sc_hd__buf_4 fanout475 (.A(net484),
    .X(net475));
 sky130_fd_sc_hd__buf_2 fanout476 (.A(net478),
    .X(net476));
 sky130_fd_sc_hd__clkbuf_2 fanout477 (.A(net478),
    .X(net477));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout478 (.A(net479),
    .X(net478));
 sky130_fd_sc_hd__buf_2 fanout479 (.A(net484),
    .X(net479));
 sky130_fd_sc_hd__buf_2 fanout480 (.A(net483),
    .X(net480));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout481 (.A(net483),
    .X(net481));
 sky130_fd_sc_hd__buf_2 fanout482 (.A(net483),
    .X(net482));
 sky130_fd_sc_hd__buf_2 fanout483 (.A(net484),
    .X(net483));
 sky130_fd_sc_hd__buf_4 fanout484 (.A(net507),
    .X(net484));
 sky130_fd_sc_hd__buf_4 fanout485 (.A(net493),
    .X(net485));
 sky130_fd_sc_hd__clkbuf_4 fanout486 (.A(net489),
    .X(net486));
 sky130_fd_sc_hd__buf_2 fanout487 (.A(net488),
    .X(net487));
 sky130_fd_sc_hd__clkbuf_2 fanout488 (.A(net489),
    .X(net488));
 sky130_fd_sc_hd__clkbuf_2 fanout489 (.A(net493),
    .X(net489));
 sky130_fd_sc_hd__buf_2 fanout490 (.A(net492),
    .X(net490));
 sky130_fd_sc_hd__buf_2 fanout491 (.A(net492),
    .X(net491));
 sky130_fd_sc_hd__clkbuf_4 fanout492 (.A(net493),
    .X(net492));
 sky130_fd_sc_hd__buf_4 fanout493 (.A(net508),
    .X(net493));
 sky130_fd_sc_hd__clkbuf_4 fanout494 (.A(net496),
    .X(net494));
 sky130_fd_sc_hd__clkbuf_2 fanout495 (.A(net496),
    .X(net495));
 sky130_fd_sc_hd__buf_2 fanout496 (.A(net506),
    .X(net496));
 sky130_fd_sc_hd__clkbuf_4 fanout497 (.A(net500),
    .X(net497));
 sky130_fd_sc_hd__buf_2 fanout498 (.A(net500),
    .X(net498));
 sky130_fd_sc_hd__clkbuf_2 fanout499 (.A(net500),
    .X(net499));
 sky130_fd_sc_hd__buf_2 fanout500 (.A(net506),
    .X(net500));
 sky130_fd_sc_hd__buf_2 fanout501 (.A(net505),
    .X(net501));
 sky130_fd_sc_hd__clkbuf_2 fanout502 (.A(net505),
    .X(net502));
 sky130_fd_sc_hd__clkbuf_4 fanout503 (.A(net505),
    .X(net503));
 sky130_fd_sc_hd__buf_2 fanout504 (.A(net505),
    .X(net504));
 sky130_fd_sc_hd__buf_2 fanout505 (.A(net506),
    .X(net505));
 sky130_fd_sc_hd__buf_4 fanout506 (.A(net508),
    .X(net506));
 sky130_fd_sc_hd__buf_6 fanout507 (.A(net46),
    .X(net507));
 sky130_fd_sc_hd__buf_4 wire508 (.A(net507),
    .X(net508));
 sky130_fd_sc_hd__conb_1 _7077__509 (.HI(net509));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_1_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_2_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_3_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_4_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_5_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_6_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_7_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_8_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_9_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_10_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_11_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_12_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_14_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_15_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_16_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_18_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_19_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_20_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_21_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_23_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_24_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_25_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_26_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_27_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_28_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_29_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_30_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_31_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_32_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_33_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_34_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_35_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_38_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_39_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_40_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_41_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_42_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_45_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_46_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_47_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_48_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_49_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_50_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_55_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_55_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_56_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_57_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_57_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_58_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_58_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_59_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_59_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_60_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_60_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_61_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_61_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_0_0_clk (.A(clknet_0_clk),
    .X(clknet_2_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_1_0_clk (.A(clknet_0_clk),
    .X(clknet_2_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_2_0_clk (.A(clknet_0_clk),
    .X(clknet_2_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_3_0_clk (.A(clknet_0_clk),
    .X(clknet_2_3_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload0 (.A(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload1 (.A(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__inv_8 clkload2 (.A(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload3 (.A(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload4 (.A(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload5 (.A(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload6 (.A(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload7 (.A(clknet_leaf_59_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload8 (.A(clknet_leaf_60_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload9 (.A(clknet_leaf_61_clk));
 sky130_fd_sc_hd__inv_6 clkload10 (.A(clknet_leaf_3_clk));
 sky130_fd_sc_hd__inv_8 clkload11 (.A(clknet_leaf_4_clk));
 sky130_fd_sc_hd__inv_6 clkload12 (.A(clknet_leaf_5_clk));
 sky130_fd_sc_hd__inv_8 clkload13 (.A(clknet_leaf_6_clk));
 sky130_fd_sc_hd__inv_8 clkload14 (.A(clknet_leaf_57_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload15 (.A(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload16 (.A(clknet_leaf_14_clk));
 sky130_fd_sc_hd__bufinv_16 clkload17 (.A(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkinv_2 clkload18 (.A(clknet_leaf_16_clk));
 sky130_fd_sc_hd__bufinv_16 clkload19 (.A(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload20 (.A(clknet_leaf_7_clk));
 sky130_fd_sc_hd__bufinv_16 clkload21 (.A(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload22 (.A(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload23 (.A(clknet_leaf_21_clk));
 sky130_fd_sc_hd__bufinv_16 clkload24 (.A(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkinv_2 clkload25 (.A(clknet_leaf_55_clk));
 sky130_fd_sc_hd__clkinv_2 clkload26 (.A(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkinv_2 clkload27 (.A(clknet_leaf_58_clk));
 sky130_fd_sc_hd__clkinv_2 clkload28 (.A(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload29 (.A(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload30 (.A(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload31 (.A(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkinv_2 clkload32 (.A(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload33 (.A(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkinv_2 clkload34 (.A(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload35 (.A(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkinv_2 clkload36 (.A(clknet_leaf_25_clk));
 sky130_fd_sc_hd__bufinv_16 clkload37 (.A(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkinv_2 clkload38 (.A(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload39 (.A(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkinv_2 clkload40 (.A(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload41 (.A(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkinv_2 clkload42 (.A(clknet_leaf_32_clk));
 sky130_fd_sc_hd__bufinv_16 clkload43 (.A(clknet_leaf_33_clk));
 sky130_fd_sc_hd__bufinv_16 clkload44 (.A(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkinv_2 clkload45 (.A(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(adc_data[3]),
    .X(net510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(net6),
    .X(net511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(adc_data[5]),
    .X(net512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(net8),
    .X(net513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(adc_data[11]),
    .X(net514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(net3),
    .X(net515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(adc_data[2]),
    .X(net516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(net5),
    .X(net517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(adc_data[1]),
    .X(net518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(net4),
    .X(net519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(adc_data[4]),
    .X(net520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(net7),
    .X(net521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(adc_data[0]),
    .X(net522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(net1),
    .X(net523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(adc_data[8]),
    .X(net524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(net11),
    .X(net525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(adc_data[7]),
    .X(net526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(net10),
    .X(net527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(adc_data[9]),
    .X(net528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(net964),
    .X(net529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(adc_valid),
    .X(net530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(net13),
    .X(net531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(_0793_),
    .X(net532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(adc_data[10]),
    .X(net533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(phase_increment[0]),
    .X(net534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(_1131_),
    .X(net535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(_0036_),
    .X(net536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(phase_increment[2]),
    .X(net537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(_1144_),
    .X(net538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(_1145_),
    .X(net539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(_0050_),
    .X(net540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(phase_increment[22]),
    .X(net541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(_1253_),
    .X(net542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(_0040_),
    .X(net543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(net812),
    .X(net544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(phase_increment[1]),
    .X(net545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(_1134_),
    .X(net546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(_1140_),
    .X(net547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(_0047_),
    .X(net548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(phase_increment[28]),
    .X(net549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(_1284_),
    .X(net550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(_0045_),
    .X(net551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(phase_increment[21]),
    .X(net552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(_1239_),
    .X(net553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(_0038_),
    .X(net554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(phase_increment[5]),
    .X(net555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(_1152_),
    .X(net556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(_1160_),
    .X(net557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(_0053_),
    .X(net558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(phase_increment[4]),
    .X(net559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(_1148_),
    .X(net560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(_1154_),
    .X(net561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(_0052_),
    .X(net562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(phase_increment[8]),
    .X(net563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(_1166_),
    .X(net564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(_0055_),
    .X(net565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(phase_increment[16]),
    .X(net566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(_1208_),
    .X(net567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(_1217_),
    .X(net568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(_0033_),
    .X(net569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(phase_increment[3]),
    .X(net570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(_1142_),
    .X(net571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(_1150_),
    .X(net572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(_0051_),
    .X(net573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(phase_increment[25]),
    .X(net574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(_0042_),
    .X(net575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(net813),
    .X(net576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(phase_increment[11]),
    .X(net577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(_1180_),
    .X(net578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(_0027_),
    .X(net579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(net815),
    .X(net580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(net814),
    .X(net581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(net818),
    .X(net582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(net822),
    .X(net583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(net816),
    .X(net584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(net819),
    .X(net585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(net817),
    .X(net586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(net833),
    .X(net587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(net835),
    .X(net588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(net824),
    .X(net589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(net826),
    .X(net590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(net839),
    .X(net591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(net834),
    .X(net592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(phase_increment[14]),
    .X(net593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(_1206_),
    .X(net594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(_0031_),
    .X(net595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(net829),
    .X(net596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(net830),
    .X(net597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(net843),
    .X(net598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(net825),
    .X(net599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(net836),
    .X(net600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(net838),
    .X(net601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(net828),
    .X(net602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(net850),
    .X(net603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(net837),
    .X(net604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(net844),
    .X(net605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(net827),
    .X(net606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(net820),
    .X(net607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(net821),
    .X(net608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(net855),
    .X(net609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(net854),
    .X(net610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(net823),
    .X(net611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(net857),
    .X(net612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(net845),
    .X(net613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(net873),
    .X(net614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(net831),
    .X(net615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(net842),
    .X(net616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(net861),
    .X(net617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(net849),
    .X(net618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(net832),
    .X(net619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(net868),
    .X(net620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(net840),
    .X(net621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(net856),
    .X(net622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(net841),
    .X(net623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(net874),
    .X(net624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(net871),
    .X(net625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(net877),
    .X(net626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(net867),
    .X(net627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(phase_increment[27]),
    .X(net628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(_0044_),
    .X(net629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(net859),
    .X(net630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(net851),
    .X(net631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(net853),
    .X(net632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(phase_increment[9]),
    .X(net633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(_1169_),
    .X(net634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(_1170_),
    .X(net635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(_0056_),
    .X(net636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(net847),
    .X(net637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(net882),
    .X(net638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(net863),
    .X(net639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(net879),
    .X(net640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(net848),
    .X(net641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(net846),
    .X(net642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(net875),
    .X(net643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(net888),
    .X(net644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(net889),
    .X(net645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(net860),
    .X(net646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(net852),
    .X(net647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(net870),
    .X(net648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(net887),
    .X(net649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(net864),
    .X(net650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(net869),
    .X(net651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(net883),
    .X(net652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(net858),
    .X(net653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(net880),
    .X(net654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(net878),
    .X(net655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(net862),
    .X(net656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(net885),
    .X(net657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(net865),
    .X(net658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(net872),
    .X(net659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(net866),
    .X(net660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(net884),
    .X(net661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(net876),
    .X(net662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(net896),
    .X(net663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(net893),
    .X(net664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(net881),
    .X(net665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(net890),
    .X(net666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(net886),
    .X(net667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(net891),
    .X(net668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(net892),
    .X(net669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(net894),
    .X(net670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(net895),
    .X(net671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(net897),
    .X(net672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(phase_increment[7]),
    .X(net673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(_1162_),
    .X(net674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(_1163_),
    .X(net675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(_0054_),
    .X(net676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(net899),
    .X(net677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(net898),
    .X(net678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(phase_increment[20]),
    .X(net679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(_1232_),
    .X(net680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(_0037_),
    .X(net681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(net900),
    .X(net682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(net901),
    .X(net683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(net902),
    .X(net684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(net930),
    .X(net685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(net927),
    .X(net686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(phase_increment[19]),
    .X(net687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(_1227_),
    .X(net688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(_1230_),
    .X(net689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(_0035_),
    .X(net690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(net924),
    .X(net691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(net925),
    .X(net692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(\mixer_q.nco_data[8] ),
    .X(net693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(net931),
    .X(net694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(phase_increment[13]),
    .X(net695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(_1192_),
    .X(net696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(_0029_),
    .X(net697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(\mixer_q.nco_data[10] ),
    .X(net698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(\mixer_q.nco_data[5] ),
    .X(net699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(net921),
    .X(net700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(net934),
    .X(net701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(net912),
    .X(net702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(net913),
    .X(net703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(net928),
    .X(net704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(phase_increment[15]),
    .X(net705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(_1211_),
    .X(net706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(_1213_),
    .X(net707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(_1214_),
    .X(net708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(_0032_),
    .X(net709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(net915),
    .X(net710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(net929),
    .X(net711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(net922),
    .X(net712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(phase_increment[30]),
    .X(net713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(_1291_),
    .X(net714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(_0048_),
    .X(net715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(net926),
    .X(net716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(net923),
    .X(net717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(net920),
    .X(net718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(net936),
    .X(net719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(phase_increment[24]),
    .X(net720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(_0041_),
    .X(net721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(net969),
    .X(net722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(phase_increment[10]),
    .X(net723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(_1176_),
    .X(net724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(_1177_),
    .X(net725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(_0026_),
    .X(net726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(phase_increment[12]),
    .X(net727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(_1190_),
    .X(net728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(_1191_),
    .X(net729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(_0028_),
    .X(net730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(\nco_inst.phase_accum[0] ),
    .X(net731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(net977),
    .X(net732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(\mixer_q.product[20] ),
    .X(net733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(\mixer_q.product[19] ),
    .X(net734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(\nco_inst.phase_accum[14] ),
    .X(net735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(_1199_),
    .X(net736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(_0030_),
    .X(net737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(\mixer_q.product[21] ),
    .X(net738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(\mixer_i.valid_stage2 ),
    .X(net739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(net967),
    .X(net740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(phase_increment[29]),
    .X(net741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(_0046_),
    .X(net742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(\nco_inst.phase_accum[21] ),
    .X(net743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(_1246_),
    .X(net744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(_1247_),
    .X(net745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(_0039_),
    .X(net746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(net970),
    .X(net747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(net968),
    .X(net748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(net971),
    .X(net749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(net932),
    .X(net750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(net975),
    .X(net751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(net933),
    .X(net752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(net953),
    .X(net753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(net935),
    .X(net754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(net958),
    .X(net755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(net954),
    .X(net756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(net962),
    .X(net757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(net942),
    .X(net758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(net960),
    .X(net759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(net956),
    .X(net760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(net943),
    .X(net761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(\mixer_i.nco_data[1] ),
    .X(net762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold254 (.A(net957),
    .X(net763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(net959),
    .X(net764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold256 (.A(net952),
    .X(net765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(net945),
    .X(net766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold258 (.A(net980),
    .X(net767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold259 (.A(net963),
    .X(net768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(net972),
    .X(net769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold261 (.A(net976),
    .X(net770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(net66),
    .X(net771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold263 (.A(net938),
    .X(net772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(net973),
    .X(net773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(net47),
    .X(net774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold266 (.A(phase_increment[17]),
    .X(net775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold267 (.A(_1220_),
    .X(net776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold268 (.A(_1225_),
    .X(net777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(_1226_),
    .X(net778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold270 (.A(net51),
    .X(net779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(net974),
    .X(net780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold272 (.A(net939),
    .X(net781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(net978),
    .X(net782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold274 (.A(net64),
    .X(net783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(net979),
    .X(net784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold276 (.A(net937),
    .X(net785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(\nco_inst.lut_addr_sin[7] ),
    .X(net786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(_1000_),
    .X(net787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(net947),
    .X(net788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(net69),
    .X(net789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(net944),
    .X(net790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(net961),
    .X(net791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold283 (.A(net946),
    .X(net792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold284 (.A(net950),
    .X(net793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold285 (.A(phase_increment[31]),
    .X(net794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold286 (.A(_1299_),
    .X(net795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(net80),
    .X(net796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold288 (.A(\mixer_i.nco_data[0] ),
    .X(net797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold289 (.A(net951),
    .X(net798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold290 (.A(net61),
    .X(net799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold291 (.A(net955),
    .X(net800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold292 (.A(\nco_inst.lut_addr_sin[6] ),
    .X(net801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold293 (.A(phase_increment[26]),
    .X(net802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold294 (.A(_1272_),
    .X(net803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold295 (.A(net965),
    .X(net804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold296 (.A(net49),
    .X(net805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold297 (.A(net83),
    .X(net806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold298 (.A(\mixer_i.nco_data[2] ),
    .X(net807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold299 (.A(net62),
    .X(net808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold300 (.A(\mixer_q.product[22] ),
    .X(net809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold301 (.A(\mixer_q.product[23] ),
    .X(net810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold302 (.A(\mixer_i.valid_stage1 ),
    .X(net811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold303 (.A(\mixer_q.product[17] ),
    .X(net812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold304 (.A(\mixer_q.product_delayed[9] ),
    .X(net813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold305 (.A(\mixer_i.product[5] ),
    .X(net814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold306 (.A(\mixer_i.product[16] ),
    .X(net815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold307 (.A(\mixer_i.product[18] ),
    .X(net816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold308 (.A(\mixer_i.product[13] ),
    .X(net817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold309 (.A(\mixer_i.nco_data[5] ),
    .X(net818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold310 (.A(\mixer_i.product[12] ),
    .X(net819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold311 (.A(\mixer_i.product_delayed[12] ),
    .X(net820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold312 (.A(\mixer_i.product[17] ),
    .X(net821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold313 (.A(\mixer_q.nco_data[2] ),
    .X(net822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold314 (.A(\mixer_i.product_delayed[3] ),
    .X(net823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold315 (.A(\mixer_i.product_delayed[8] ),
    .X(net824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold316 (.A(\mixer_i.product[11] ),
    .X(net825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold317 (.A(\mixer_i.product_delayed[7] ),
    .X(net826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold318 (.A(\mixer_i.product[8] ),
    .X(net827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold319 (.A(\mixer_i.product[7] ),
    .X(net828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold320 (.A(\mixer_i.product_delayed[15] ),
    .X(net829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold321 (.A(\mixer_i.product_delayed[13] ),
    .X(net830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold322 (.A(\mixer_i.product_delayed[21] ),
    .X(net831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold323 (.A(\mixer_i.product_delayed[9] ),
    .X(net832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold324 (.A(\mixer_q.nco_data[1] ),
    .X(net833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold325 (.A(\mixer_q.product[4] ),
    .X(net834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold326 (.A(\mixer_q.nco_data[3] ),
    .X(net835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold327 (.A(\mixer_q.product_delayed[22] ),
    .X(net836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold328 (.A(\mixer_i.product_delayed[0] ),
    .X(net837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold329 (.A(\mixer_i.product_delayed[6] ),
    .X(net838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold330 (.A(\mixer_i.product[6] ),
    .X(net839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold331 (.A(\mixer_i.product_delayed[2] ),
    .X(net840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold332 (.A(\mixer_i.product[3] ),
    .X(net841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold333 (.A(\mixer_q.product_delayed[19] ),
    .X(net842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold334 (.A(\mixer_q.nco_data[0] ),
    .X(net843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold335 (.A(\mixer_i.nco_data[3] ),
    .X(net844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold336 (.A(\mixer_q.product_delayed[21] ),
    .X(net845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold337 (.A(\mixer_i.product_delayed[20] ),
    .X(net846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold338 (.A(\mixer_q.product_delayed[23] ),
    .X(net847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold339 (.A(\mixer_i.valid_stage2_delayed ),
    .X(net848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold340 (.A(\mixer_q.product[16] ),
    .X(net849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold341 (.A(\mixer_q.product_delayed[10] ),
    .X(net850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold342 (.A(\mixer_i.product[14] ),
    .X(net851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold343 (.A(\mixer_i.product[1] ),
    .X(net852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold344 (.A(\mixer_q.product[6] ),
    .X(net853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold345 (.A(\mixer_q.product[13] ),
    .X(net854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold346 (.A(\mixer_q.product_delayed[5] ),
    .X(net855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold347 (.A(\mixer_i.product[15] ),
    .X(net856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold348 (.A(\mixer_q.product[11] ),
    .X(net857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold349 (.A(\mixer_q.product_delayed[1] ),
    .X(net858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold350 (.A(\mixer_i.product[4] ),
    .X(net859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold351 (.A(\mixer_q.product[2] ),
    .X(net860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold352 (.A(\mixer_q.product_delayed[7] ),
    .X(net861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold353 (.A(\mixer_i.product_delayed[16] ),
    .X(net862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold354 (.A(\mixer_i.product[10] ),
    .X(net863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold355 (.A(\mixer_q.product_delayed[3] ),
    .X(net864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold356 (.A(\mixer_i.product[0] ),
    .X(net865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold357 (.A(\mixer_i.product_delayed[23] ),
    .X(net866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold358 (.A(\mixer_q.product_delayed[11] ),
    .X(net867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold359 (.A(\mixer_q.product_delayed[6] ),
    .X(net868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold360 (.A(\mixer_q.product_delayed[12] ),
    .X(net869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold361 (.A(\mixer_i.product[23] ),
    .X(net870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold362 (.A(\mixer_q.product[10] ),
    .X(net871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold363 (.A(\mixer_i.product_delayed[22] ),
    .X(net872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold364 (.A(\mixer_q.product_delayed[16] ),
    .X(net873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold365 (.A(\mixer_q.product[15] ),
    .X(net874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold366 (.A(\mixer_q.nco_data[4] ),
    .X(net875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold367 (.A(\mixer_i.product_delayed[11] ),
    .X(net876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold368 (.A(\mixer_q.product_delayed[15] ),
    .X(net877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold369 (.A(\mixer_q.product_delayed[8] ),
    .X(net878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold370 (.A(\mixer_q.product[8] ),
    .X(net879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold371 (.A(\mixer_q.product[3] ),
    .X(net880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold372 (.A(\mixer_i.product_delayed[5] ),
    .X(net881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold373 (.A(\mixer_q.product[5] ),
    .X(net882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold374 (.A(\mixer_i.nco_data[4] ),
    .X(net883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold375 (.A(\mixer_q.product_delayed[4] ),
    .X(net884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold376 (.A(\mixer_q.nco_data[7] ),
    .X(net885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold377 (.A(\mixer_q.product_delayed[20] ),
    .X(net886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold378 (.A(\mixer_q.product_delayed[13] ),
    .X(net887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold379 (.A(\mixer_q.product[14] ),
    .X(net888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold380 (.A(\mixer_q.product_delayed[14] ),
    .X(net889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold381 (.A(\mixer_q.product[12] ),
    .X(net890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold382 (.A(\mixer_i.nco_data[9] ),
    .X(net891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold383 (.A(\mixer_i.product_delayed[19] ),
    .X(net892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold384 (.A(\mixer_q.product[7] ),
    .X(net893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold385 (.A(\mixer_i.product[2] ),
    .X(net894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold386 (.A(\mixer_q.product[0] ),
    .X(net895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold387 (.A(\mixer_q.nco_data[6] ),
    .X(net896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold388 (.A(\mixer_q.product_delayed[17] ),
    .X(net897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold389 (.A(\mixer_i.product_delayed[4] ),
    .X(net898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold390 (.A(\mixer_q.nco_data[9] ),
    .X(net899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold391 (.A(\mixer_i.product[9] ),
    .X(net900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold392 (.A(\mixer_q.product_delayed[18] ),
    .X(net901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold393 (.A(\mixer_i.product_delayed[14] ),
    .X(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_0062_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_0062_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_0073_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_0074_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_0074_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_0133_));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_0221_));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_0365_));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_0385_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(_0385_));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(_0395_));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(_0802_));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(_0802_));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(_0818_));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(_0912_));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(_0946_));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(_0965_));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(_1166_));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(_1214_));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(_1329_));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(_1329_));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(_1329_));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(_1782_));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(_1810_));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(_1869_));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(_1933_));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(_1985_));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(_2218_));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(_2848_));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(_2973_));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(_2973_));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(_3058_));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(_3125_));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(_3125_));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(_3134_));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(_3176_));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(_3176_));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(_3178_));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(_3178_));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(_3178_));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(_3182_));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(_3355_));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(_3355_));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(_3394_));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(_3441_));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(_3455_));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(_3475_));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(_3475_));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(\mixer_i.adc_reg[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(\mixer_i.adc_reg[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(\mixer_i.adc_reg[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(\mixer_i.adc_reg[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(\mixer_i.nco_reg[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(\mixer_i.nco_reg[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(\mixer_i.valid_stage1 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(\mixer_q.nco_reg[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(\mixer_q.nco_reg[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(\mixer_q.nco_reg[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(\mixer_q.nco_reg[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(\mixer_q.nco_reg[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(\mixer_q.nco_reg[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(\mixer_q.nco_reg[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(\mixer_q.product[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(\mixer_q.product[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_73 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_74 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_75 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_76 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_77 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_78 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_79 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_80 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_81 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_82 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_83 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_84 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_85 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_86 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA_87 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_88 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_89 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_90 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_91 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_92 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_93 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_94 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_95 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_96 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_97 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_98 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA_99 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_100 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_101 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_102 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA_103 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA_104 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_105 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_106 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_107 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_108 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_109 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_110 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA_111 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA_112 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_113 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_114 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_115 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_116 (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA_117 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA_118 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA_119 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_120 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_121 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_122 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_123 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_124 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_125 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA_126 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_127 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_128 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_129 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_130 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_131 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA_132 (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA_133 (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA_134 (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA_135 (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA_136 (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA_137 (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA_138 (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA_139 (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA_140 (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 ANTENNA_141 (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 ANTENNA_142 (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 ANTENNA_143 (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 ANTENNA_144 (.DIODE(net507));
 sky130_fd_sc_hd__diode_2 ANTENNA_145 (.DIODE(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_146 (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_147 (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA_148 (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_149 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_150 (.DIODE(_0509_));
 sky130_fd_sc_hd__diode_2 ANTENNA_151 (.DIODE(_0509_));
 sky130_fd_sc_hd__diode_2 ANTENNA_152 (.DIODE(_0737_));
 sky130_fd_sc_hd__diode_2 ANTENNA_153 (.DIODE(_0737_));
 sky130_fd_sc_hd__diode_2 ANTENNA_154 (.DIODE(_0912_));
 sky130_fd_sc_hd__diode_2 ANTENNA_155 (.DIODE(_1329_));
 sky130_fd_sc_hd__diode_2 ANTENNA_156 (.DIODE(_1394_));
 sky130_fd_sc_hd__diode_2 ANTENNA_157 (.DIODE(_1407_));
 sky130_fd_sc_hd__diode_2 ANTENNA_158 (.DIODE(_2093_));
 sky130_fd_sc_hd__diode_2 ANTENNA_159 (.DIODE(_2794_));
 sky130_fd_sc_hd__diode_2 ANTENNA_160 (.DIODE(_3134_));
 sky130_fd_sc_hd__diode_2 ANTENNA_161 (.DIODE(_3179_));
 sky130_fd_sc_hd__diode_2 ANTENNA_162 (.DIODE(_3228_));
 sky130_fd_sc_hd__diode_2 ANTENNA_163 (.DIODE(_3441_));
 sky130_fd_sc_hd__diode_2 ANTENNA_164 (.DIODE(\mixer_i.adc_reg[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_165 (.DIODE(\mixer_i.adc_reg[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_166 (.DIODE(\mixer_i.valid_stage2 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_167 (.DIODE(\mixer_q.nco_reg[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_168 (.DIODE(\nco_inst.cosine_lut.addr[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_169 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_170 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_171 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_172 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_173 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_174 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_175 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_176 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_177 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_178 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_179 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_180 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_181 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA_182 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA_183 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA_184 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA_185 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA_186 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_187 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_188 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA_189 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA_190 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_191 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_192 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_193 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_194 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_195 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_196 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_197 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_198 (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA_199 (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA_200 (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA_201 (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_202 (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_203 (.DIODE(_0509_));
 sky130_fd_sc_hd__diode_2 ANTENNA_204 (.DIODE(_0810_));
 sky130_fd_sc_hd__diode_2 ANTENNA_205 (.DIODE(_0905_));
 sky130_fd_sc_hd__diode_2 ANTENNA_206 (.DIODE(_1407_));
 sky130_fd_sc_hd__diode_2 ANTENNA_207 (.DIODE(_3058_));
 sky130_fd_sc_hd__diode_2 ANTENNA_208 (.DIODE(_3134_));
 sky130_fd_sc_hd__diode_2 ANTENNA_209 (.DIODE(\mixer_i.adc_reg[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_210 (.DIODE(\nco_inst.cosine_lut.addr[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_211 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_212 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA_213 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_214 (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA_215 (.DIODE(_0057_));
 sky130_fd_sc_hd__diode_2 ANTENNA_216 (.DIODE(_0057_));
 sky130_fd_sc_hd__diode_2 ANTENNA_217 (.DIODE(_0810_));
 sky130_fd_sc_hd__diode_2 ANTENNA_218 (.DIODE(_3058_));
 sky130_fd_sc_hd__diode_2 ANTENNA_219 (.DIODE(_3058_));
 sky130_fd_sc_hd__diode_2 ANTENNA_220 (.DIODE(_0810_));
 sky130_fd_sc_hd__diode_2 ANTENNA_221 (.DIODE(net376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold395 (.A(net174),
    .X(net904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold397 (.A(net698),
    .X(net906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold398 (.A(\mixer_i.nco_reg[2] ),
    .X(net907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold399 (.A(_2817_),
    .X(net908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold400 (.A(_2865_),
    .X(net909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold401 (.A(_2875_),
    .X(net910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold402 (.A(_0100_),
    .X(net911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold403 (.A(\mixer_q.product[9] ),
    .X(net912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold404 (.A(\mixer_q.nco_data[11] ),
    .X(net913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold405 (.A(\nco_inst.cosine_lut.addr[1] ),
    .X(net914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold406 (.A(\mixer_i.nco_data[8] ),
    .X(net915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold408 (.A(net699),
    .X(net917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold410 (.A(net693),
    .X(net919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold411 (.A(\mixer_i.nco_data[10] ),
    .X(net920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold412 (.A(\mixer_q.product_delayed[2] ),
    .X(net921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold413 (.A(\mixer_i.nco_data[6] ),
    .X(net922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold414 (.A(\mixer_i.nco_data[7] ),
    .X(net923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold415 (.A(\mixer_i.product[19] ),
    .X(net924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold416 (.A(\mixer_q.product_delayed[0] ),
    .X(net925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold417 (.A(\mixer_i.nco_data[11] ),
    .X(net926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold418 (.A(\mixer_i.product_delayed[18] ),
    .X(net927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold419 (.A(\mixer_i.product[22] ),
    .X(net928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold420 (.A(\mixer_q.product[1] ),
    .X(net929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold421 (.A(\mixer_i.product_delayed[10] ),
    .X(net930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold422 (.A(\mixer_i.product_delayed[17] ),
    .X(net931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold423 (.A(net50),
    .X(net932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold424 (.A(net52),
    .X(net933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold425 (.A(\mixer_i.product_delayed[1] ),
    .X(net934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold426 (.A(net95),
    .X(net935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold427 (.A(\mixer_i.product[20] ),
    .X(net936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold428 (.A(net91),
    .X(net937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold429 (.A(net82),
    .X(net938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold430 (.A(net87),
    .X(net939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold431 (.A(\mixer_i.nco_reg[1] ),
    .X(net940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold432 (.A(_2827_),
    .X(net941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold433 (.A(net54),
    .X(net942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold434 (.A(net55),
    .X(net943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold435 (.A(net92),
    .X(net944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold436 (.A(net56),
    .X(net945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold437 (.A(net94),
    .X(net946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold438 (.A(net93),
    .X(net947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold440 (.A(net779),
    .X(net949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold441 (.A(net90),
    .X(net950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold442 (.A(net89),
    .X(net951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold443 (.A(net57),
    .X(net952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold444 (.A(net72),
    .X(net953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold445 (.A(net78),
    .X(net954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold446 (.A(net88),
    .X(net955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold447 (.A(net73),
    .X(net956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold448 (.A(net74),
    .X(net957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold449 (.A(net77),
    .X(net958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold450 (.A(net75),
    .X(net959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold451 (.A(net59),
    .X(net960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold452 (.A(net53),
    .X(net961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold453 (.A(net76),
    .X(net962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold454 (.A(net60),
    .X(net963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold455 (.A(adc_data[6]),
    .X(net964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold456 (.A(net71),
    .X(net965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold457 (.A(\nco_inst.cosine_lut.addr[5] ),
    .X(net966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold458 (.A(net84),
    .X(net967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold459 (.A(net81),
    .X(net968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold460 (.A(\mixer_i.product[21] ),
    .X(net969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold461 (.A(net79),
    .X(net970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold462 (.A(net85),
    .X(net971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold463 (.A(net48),
    .X(net972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold464 (.A(net68),
    .X(net973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold465 (.A(net67),
    .X(net974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold466 (.A(net86),
    .X(net975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold467 (.A(net65),
    .X(net976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold468 (.A(\mixer_q.product[18] ),
    .X(net977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold469 (.A(net70),
    .X(net978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold470 (.A(net58),
    .X(net979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold471 (.A(net63),
    .X(net980));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1329 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1341 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_1349 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1343 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_1345 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1353 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1329 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1337 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1359 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1315 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1337 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1354 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1362 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1269 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1277 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1280 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1277 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1298 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1325 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1337 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_1349 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1257 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1269 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1275 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1278 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1309 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1321 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1329 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1339 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1273 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1315 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1352 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1363 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1296 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1308 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_1361 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1287 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1297 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1305 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_1341 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1351 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1261 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1310 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1337 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1289 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1320 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1332 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1363 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1281 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1293 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1305 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_1361 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1265 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_1277 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1363 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1361 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1361 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1297 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1309 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1321 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1333 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1270 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1282 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1310 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1322 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1334 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1342 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1351 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1261 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_1283 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1302 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1317 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1352 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1363 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1217 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1235 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1277 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_1361 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1297 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1309 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1321 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1333 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_1361 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1363 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1329 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1341 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_1349 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_18 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1329 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1075 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1111 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1301 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1333 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1064 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1281 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1299 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1303 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_1361 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_635 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1207 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1265 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1277 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1321 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1333 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1173 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1203 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_1210 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1220 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1228 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1281 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1293 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1305 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_1361 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_995 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1098 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1287 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1311 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1320 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1332 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1164 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1184 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1241 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1273 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1298 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1310 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1175 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1187 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1256 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_1264 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1343 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1351 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1189 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1229 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1329 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1333 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1362 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1363 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1102 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1173 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1244 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1273 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1285 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1293 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1315 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1337 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1349 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_1361 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1138 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1203 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1215 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1240 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1249 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1265 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1286 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1324 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1336 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_875 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_878 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_886 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_904 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1129 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1202 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_1209 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1238 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1273 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_873 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_929 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1036 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1128 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1135 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1183 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1195 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1207 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1219 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1266 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1278 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1363 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_955 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1055 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1067 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1218 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1222 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1234 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_1361 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_929 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1038 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1110 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1114 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1131 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1141 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1190 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1214 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1103 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1152 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1259 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1268 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1274 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1295 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1317 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_1341 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1360 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_870 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_882 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1189 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1201 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1287 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1295 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1312 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_1334 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1342 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1351 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_6 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_970 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_974 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1008 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1012 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1120 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1202 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1243 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1265 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1277 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_917 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1192 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_1204 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1269 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1281 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_888 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_908 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_936 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_958 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_998 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1010 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1018 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1030 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1047 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1171 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1259 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1261 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1269 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1278 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1286 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1312 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1337 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_1257 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1271 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1283 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1287 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1340 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_1061 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_1069 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1078 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1086 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1135 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1223 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1235 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1285 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_1297 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_1305 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1337 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_868 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_917 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_927 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1096 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1119 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1197 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1266 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1278 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1301 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1323 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1335 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1185 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1196 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1223 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1237 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1259 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1265 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1341 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_1353 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1194 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1206 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1230 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1239 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1263 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1343 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1345 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_1353 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1011 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_1361 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_870 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_918 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_936 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_970 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1038 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1060 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1087 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_1098 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_1129 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_1155 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1309 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1321 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1333 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_1341 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1351 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1116 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1122 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1128 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1341 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_873 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1056 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1270 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1282 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1363 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_938 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_974 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1008 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1032 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1067 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1225 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1239 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_1361 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1038 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_1050 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1085 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1098 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1243 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1266 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1278 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1286 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1305 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1319 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1331 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1363 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_945 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1044 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1080 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_1086 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1259 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1290 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_1361 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1098 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1266 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1278 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1332 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_880 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1113 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1229 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1261 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1310 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1317 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1325 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1355 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_900 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_926 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_938 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1287 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1296 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1309 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1321 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_1333 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1125 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1244 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1285 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1297 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1329 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1341 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_1349 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1289 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1324 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1336 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1363 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_844 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_882 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_952 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1102 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1110 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_1246 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_1361 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_991 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_1309 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1332 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1153 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1222 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1234 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1317 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_1329 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1360 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1208 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1363 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1069 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1083 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1106 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_1114 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1120 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_1128 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1159 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_1171 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1315 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1317 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_1325 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1336 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1348 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_863 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_875 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1089 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1343 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_1345 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_1353 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_910 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1119 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_1313 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1339 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1124 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1200 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1225 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1293 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1305 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1329 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1341 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_1349 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1135 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_884 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1097 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1112 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1120 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1212 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1236 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_860 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1056 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1095 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_1103 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1131 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1180 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1192 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1206 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1109 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1124 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1159 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1171 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1183 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1244 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1341 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1353 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1362 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_816 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_964 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1125 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1132 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_945 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1242 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1278 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1290 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1302 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1329 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1333 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1354 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1362 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_814 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1175 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1187 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1271 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1283 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1343 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1353 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1362 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1029 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1146 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1181 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1244 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1281 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1293 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1305 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1341 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1353 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1362 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_690 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_714 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1131 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1199 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1343 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1351 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1167 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1187 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1240 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_961 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1229 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_1236 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_1361 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_749 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1026 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1038 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1253 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1265 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1280 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1363 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1004 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_1011 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1066 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1109 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1155 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1179 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1191 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_688 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1040 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_1051 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1103 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1172 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1187 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1363 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_882 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_912 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_916 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1111 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1153 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1244 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_1361 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_807 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_868 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_901 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1098 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1222 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1260 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_1272 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1363 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_857 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1223 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1235 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1259 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1265 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1270 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1296 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_1308 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_1201 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1270 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1343 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1351 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1046 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1229 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1261 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1282 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1294 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_1306 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_644 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_702 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_970 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1145 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1169 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_1183 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1199 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1255 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1267 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1363 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_886 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1047 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1059 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1162 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_1361 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_734 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1036 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1060 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1116 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_1185 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1204 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_1216 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1245 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_1257 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_1265 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1271 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1275 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_1280 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1363 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_620 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1173 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1200 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1225 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_1236 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_1244 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1261 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1325 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1337 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1349 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1355 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_536 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_940 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1197 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1258 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1263 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1287 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_1333 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_1341 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_1353 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_507 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_539 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_665 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_804 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1185 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1242 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1254 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1268 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_1276 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_1284 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1307 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1328 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1332 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_693 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1190 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1208 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1271 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1283 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1309 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1318 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1330 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1342 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1351 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_732 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_972 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1010 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1153 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1171 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1183 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1223 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1270 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1282 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1294 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1306 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1337 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1361 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_970 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_982 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1137 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1189 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1226 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_1236 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1249 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1267 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1313 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_1325 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_1333 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_1361 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_679 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_777 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_929 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_1253 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1269 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1275 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1281 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1293 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1309 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_1361 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_759 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_861 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_927 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_956 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1138 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1150 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1243 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1263 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1310 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1323 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_1335 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_808 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1091 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1100 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1229 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1247 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1285 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_1297 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_1305 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1352 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1016 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_1040 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1048 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1301 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1313 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1317 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1338 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_1345 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1353 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_988 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1000 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1012 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1050 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1107 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_1126 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_1215 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1223 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1242 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1281 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1293 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_1361 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1045 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1324 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_1336 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_1345 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_1353 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_778 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_885 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1109 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1315 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1337 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_1361 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_817 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_948 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1174 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1191 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1208 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1301 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1313 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_1325 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_1333 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_1361 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_788 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_806 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_930 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1281 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1299 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_1337 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1348 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_471 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1036 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1343 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_679 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1048 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_1084 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1112 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_1185 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1063 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1114 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1200 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1262 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_822 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_972 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1010 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1054 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1066 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1078 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1113 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1183 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_1188 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1341 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_1353 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1041 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_1056 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_1075 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1139 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_1151 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1163 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1270 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1282 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_891 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_914 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1225 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_1098 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1128 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1152 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_1164 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1343 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_1345 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_1353 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_723 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_935 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1221 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1236 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1275 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1299 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1340 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1352 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_579 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_812 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1098 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1118 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1209 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1215 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1287 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1315 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1340 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1351 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1064 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1156 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1208 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1239 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1285 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_1297 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_1305 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1337 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1349 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1355 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_690 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1118 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1170 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1221 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1255 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1267 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1322 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_1334 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1176 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_1188 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1202 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_1222 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1238 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1363 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1010 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1176 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_1188 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1240 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_901 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_919 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_917 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1017 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1055 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_1067 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1109 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1136 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1166 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1183 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_807 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_980 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_992 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1092 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1131 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1143 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_1173 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_1184 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1212 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1343 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_945 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1008 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1069 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1104 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1112 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_1124 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_539 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_944 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1343 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1351 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_539 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_833 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_842 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1152 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1261 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1273 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1299 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1303 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_946 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1063 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1098 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1287 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1296 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1326 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1338 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_827 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1066 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1070 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1097 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1102 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1110 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1122 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1159 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_1171 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_1212 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1237 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1317 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1352 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_588 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_870 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1053 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1171 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1194 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1216 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1220 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_1224 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1255 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1267 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1313 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1343 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_1361 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1001 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1059 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1124 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1152 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1164 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1168 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_1218 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_1226 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_1236 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1243 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_1252 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1295 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_1307 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1317 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1329 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1335 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_1356 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_844 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1089 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1183 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1195 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1207 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1240 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1263 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1343 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_1345 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_1353 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1050 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1086 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1120 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_1168 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1182 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1222 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1234 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1258 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1282 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1304 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1341 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1353 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1363 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_532 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_974 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_994 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1174 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1208 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1245 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_1257 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_1265 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1331 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1363 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_884 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_999 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1173 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1191 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1208 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1220 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1329 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1341 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_1349 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_532 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_966 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1036 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1119 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1181 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1363 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_959 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_994 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1091 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_1173 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1219 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1224 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_1361 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1094 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1174 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1184 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1202 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1236 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1248 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1260 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1363 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1064 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1103 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_1115 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_1123 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1146 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1199 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1281 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1293 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_1305 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_1313 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1326 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1338 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1350 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1362 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1039 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1212 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1238 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_969 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1062 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1079 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_1145 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1170 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_1182 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1190 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1235 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1285 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_1305 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_1329 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1337 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1359 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_812 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_924 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_935 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1018 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1038 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1195 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1210 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1230 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1270 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1282 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1343 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_1345 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_1353 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1091 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_1103 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1203 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1218 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1230 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_1234 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1299 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1315 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1341 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_1353 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_760 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_1141 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_1229 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1262 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_779 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_969 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1153 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1182 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_1194 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1223 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_1235 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1259 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1298 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1310 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1329 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_1341 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_1349 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1015 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1050 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1145 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1212 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1245 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_1257 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_1265 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1303 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1327 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1339 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_966 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1017 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1061 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1259 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1265 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1286 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_1361 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1072 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1183 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1195 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1207 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1287 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1297 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1320 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1332 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1363 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1153 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1178 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1215 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1227 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1239 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_1361 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_534 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_907 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_918 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1297 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1309 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1321 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_1333 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1363 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_864 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_891 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_907 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1147 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_878 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_929 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1094 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_1185 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1210 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1301 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_1313 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_1321 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_499 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1081 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1223 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1235 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1273 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1341 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_804 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_816 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1004 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1075 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1208 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1287 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1324 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_1336 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1351 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_888 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1066 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1089 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1107 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_901 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_939 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1155 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_1361 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_14 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_822 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1085 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1139 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1363 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_450 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_658 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_723 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_957 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_991 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1273 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_1285 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_1293 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_1361 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_666 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1051 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1297 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1317 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1363 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_936 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_960 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_992 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1004 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1317 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_1337 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1360 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_973 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1287 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1332 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_1345 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_1353 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_844 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_855 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_916 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_939 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_947 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_995 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1315 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1317 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1326 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1332 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_1353 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_666 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1343 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1351 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_678 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_936 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_964 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_535 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1008 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_665 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_799 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_902 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_948 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1024 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_1036 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_886 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_952 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1287 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1325 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_1334 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_609 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1315 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1321 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1330 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1352 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_703 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_807 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_946 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1026 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1038 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1343 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_1345 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_946 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_966 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1050 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1329 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_1341 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_1349 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_639 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_799 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1039 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_916 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_888 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1305 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1321 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_1333 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_819 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_982 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1019 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1039 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1343 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_1345 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_731 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1273 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1325 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1337 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1349 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1309 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1338 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_883 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_816 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1343 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_784 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_882 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_935 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1047 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1059 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1329 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_1341 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_1349 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_1040 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1001 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1008 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1051 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_532 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_994 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1051 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_791 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_964 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_957 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_963 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_995 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1054 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1066 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_946 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_962 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_823 ();
 sky130_fd_sc_hd__decap_3 FILLER_212_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_212_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_212_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1042 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1046 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_212_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_213_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_213_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_213_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_870 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_1056 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1343 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1351 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_1086 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1063 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_216_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_216_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_216_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_1004 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_1036 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1078 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1114 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_217_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1214 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1363 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1016 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_1030 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_1185 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1237 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_1361 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_219_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_219_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_219_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_219_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_907 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_1036 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_1058 ();
 sky130_fd_sc_hd__decap_3 FILLER_219_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1098 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_219_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_220_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_220_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_220_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1189 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_220_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1236 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_220_1281 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1298 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_1310 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_220_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_221_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_221_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_221_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_221_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_221_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_221_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1039 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_221_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_222_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_222_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_222_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_222_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_222_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_222_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_222_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1239 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_222_1281 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1304 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_222_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_223_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_223_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_223_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_223_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_223_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_223_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_223_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_223_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_799 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_929 ();
 sky130_fd_sc_hd__decap_3 FILLER_223_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_223_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1023 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1098 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1153 ();
 sky130_fd_sc_hd__decap_3 FILLER_223_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1320 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1332 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1351 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_224_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_224_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_224_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_224_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_224_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_224_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_224_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_224_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_224_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1285 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_1297 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1307 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1337 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1349 ();
 sky130_fd_sc_hd__decap_3 FILLER_224_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_225_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_225_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_225_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_722 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_225_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_225_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1343 ();
 sky130_fd_sc_hd__decap_3 FILLER_225_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_1117 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_1341 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1363 ();
endmodule
